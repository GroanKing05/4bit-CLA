magic
tech scmos
timestamp 1731497959
<< nwell >>
rect -22 219 12 239
rect -22 187 45 219
rect 56 202 88 235
rect 68 163 93 195
<< ntransistor >>
rect 95 222 105 224
rect 95 213 105 215
rect -11 165 -9 175
rect -1 165 1 175
rect 22 155 24 175
rect 32 155 34 175
rect 79 147 81 157
<< ptransistor >>
rect -11 193 -9 233
rect -1 193 1 233
rect 62 222 82 224
rect 62 213 82 215
rect 22 193 24 213
rect 32 193 34 213
rect 79 169 81 189
<< ndiffusion >>
rect 99 225 105 229
rect 95 224 105 225
rect 95 220 105 222
rect 99 216 105 220
rect 95 215 105 216
rect 95 212 105 213
rect 95 208 101 212
rect -16 169 -11 175
rect -12 165 -11 169
rect -9 171 -7 175
rect -3 171 -1 175
rect -9 165 -1 171
rect 1 169 6 175
rect 1 165 2 169
rect 17 159 22 175
rect 21 155 22 159
rect 24 155 32 175
rect 34 171 35 175
rect 34 155 39 171
rect 74 151 79 157
rect 78 147 79 151
rect 81 153 82 157
rect 81 147 86 153
<< pdiffusion >>
rect -16 197 -11 233
rect -12 193 -11 197
rect -9 193 -1 233
rect 1 229 2 233
rect 1 193 6 229
rect 62 225 78 229
rect 62 224 82 225
rect 62 220 82 222
rect 62 216 76 220
rect 80 216 82 220
rect 62 215 82 216
rect 21 209 22 213
rect 17 193 22 209
rect 24 197 32 213
rect 24 193 26 197
rect 30 193 32 197
rect 34 209 35 213
rect 34 193 39 209
rect 62 212 82 213
rect 66 208 82 212
rect 78 185 79 189
rect 74 169 79 185
rect 81 173 86 189
rect 81 169 82 173
<< ndcontact >>
rect 95 225 99 229
rect 95 216 99 220
rect 101 208 105 212
rect -16 165 -12 169
rect -7 171 -3 175
rect 2 165 6 169
rect 17 155 21 159
rect 35 171 39 175
rect 74 147 78 151
rect 82 153 86 157
<< pdcontact >>
rect -16 193 -12 197
rect 2 229 6 233
rect 78 225 82 229
rect 76 216 80 220
rect 17 209 21 213
rect 26 193 30 197
rect 35 209 39 213
rect 62 208 66 212
rect 74 185 78 189
rect 82 169 86 173
<< polysilicon >>
rect -11 233 -9 236
rect -1 233 1 236
rect 50 222 62 224
rect 82 222 88 224
rect 91 222 95 224
rect 105 223 112 224
rect 105 222 107 223
rect 22 213 24 217
rect 32 213 34 217
rect 111 222 112 223
rect 59 213 62 215
rect 82 213 95 215
rect 105 213 108 215
rect -11 175 -9 193
rect -1 175 1 193
rect 22 175 24 193
rect 32 175 34 193
rect 79 189 81 193
rect -11 162 -9 165
rect -1 162 1 165
rect 79 157 81 169
rect 22 151 24 155
rect 32 151 34 155
rect 79 143 81 147
<< polycontact >>
rect 51 218 55 222
rect 107 219 111 223
rect 89 209 93 213
rect -9 182 -5 186
rect 18 183 22 187
rect 1 176 5 180
rect 28 176 32 180
rect 75 158 79 162
<< metal1 >>
rect -22 240 8 243
rect 50 241 92 244
rect 3 233 6 240
rect 9 223 12 240
rect 89 237 92 241
rect 89 232 91 237
rect 89 228 92 232
rect 82 225 95 228
rect 9 220 45 223
rect 17 213 20 220
rect 35 213 39 220
rect 52 200 55 218
rect 80 217 83 220
rect 88 217 95 220
rect 51 199 55 200
rect 62 199 65 208
rect 90 203 93 209
rect 102 205 105 208
rect 108 205 111 219
rect 51 196 65 199
rect 73 196 77 199
rect 100 202 111 205
rect -16 184 -13 193
rect 9 186 12 193
rect 27 192 30 193
rect 27 189 39 192
rect -22 181 -13 184
rect -5 183 18 186
rect -16 179 -13 181
rect 36 180 39 189
rect -16 176 -4 179
rect 5 177 28 180
rect -7 175 -4 176
rect 9 173 12 177
rect 36 177 45 180
rect 36 175 39 177
rect -16 161 -13 165
rect 3 161 6 165
rect 62 162 65 196
rect 74 189 77 196
rect 100 192 103 202
rect 94 189 103 192
rect 83 162 86 169
rect 94 162 97 189
rect -22 158 14 161
rect 62 159 75 162
rect 11 150 14 158
rect 83 159 97 162
rect 83 157 86 159
rect 17 150 20 155
rect 11 147 74 150
<< m2contact >>
rect 8 240 14 245
rect 45 240 50 245
rect 83 216 88 221
rect 9 193 14 198
rect 46 195 51 200
rect 68 196 73 201
rect 9 168 14 173
<< metal2 >>
rect 35 250 72 253
rect 35 244 38 250
rect 14 241 38 244
rect 46 229 49 240
rect 10 226 50 229
rect 10 198 13 226
rect 26 215 50 218
rect 26 172 29 215
rect 47 200 50 215
rect 69 201 72 250
rect 84 221 87 237
rect 14 169 29 172
<< m123contact >>
rect 91 232 96 237
rect 89 198 94 203
<< metal3 >>
rect 90 232 91 235
rect 90 203 93 232
<< labels >>
rlabel metal1 5 241 5 242 5 vdd
rlabel metal1 -5 160 -5 160 1 gnd
rlabel metal1 23 221 23 221 5 vdd
rlabel metal1 32 148 32 148 1 gnd
rlabel metal1 6 183 17 186 1 in1
rlabel metal1 7 177 13 180 1 in2
rlabel metal2 47 226 50 229 1 in1
rlabel metal2 47 215 50 218 1 in2
rlabel metal1 -21 181 -17 183 3 p_inv
rlabel metal1 39 177 45 180 1 g_inv
rlabel metal3 90 230 90 230 7 in2
rlabel metal1 89 218 89 218 7 out
rlabel metal1 75 197 75 197 7 vdd
rlabel metal1 69 159 72 161 3 in1
rlabel metal1 85 160 85 160 1 in1_inv
<< end >>
