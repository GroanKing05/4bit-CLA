magic
tech scmos
timestamp 1731589888
<< nwell >>
rect -191 -85 -130 -53
<< ntransistor >>
rect -180 -101 -178 -91
rect -152 -102 -150 -92
rect -143 -102 -141 -92
<< ptransistor >>
rect -180 -79 -178 -59
rect -152 -79 -150 -59
rect -143 -79 -141 -59
<< ndiffusion >>
rect -185 -97 -180 -91
rect -181 -101 -180 -97
rect -178 -97 -173 -91
rect -178 -101 -177 -97
rect -157 -98 -152 -92
rect -153 -102 -152 -98
rect -150 -96 -149 -92
rect -145 -96 -143 -92
rect -150 -102 -143 -96
rect -141 -96 -140 -92
rect -141 -102 -136 -96
<< pdiffusion >>
rect -185 -75 -180 -59
rect -181 -79 -180 -75
rect -178 -63 -177 -59
rect -178 -79 -173 -63
rect -153 -63 -152 -59
rect -157 -79 -152 -63
rect -150 -73 -143 -59
rect -150 -77 -149 -73
rect -145 -77 -143 -73
rect -150 -79 -143 -77
rect -141 -75 -136 -59
rect -141 -79 -140 -75
<< ndcontact >>
rect -185 -101 -181 -97
rect -177 -101 -173 -97
rect -157 -102 -153 -98
rect -149 -96 -145 -92
rect -140 -96 -136 -92
<< pdcontact >>
rect -185 -79 -181 -75
rect -177 -63 -173 -59
rect -157 -63 -153 -59
rect -149 -77 -145 -73
rect -140 -79 -136 -75
<< polysilicon >>
rect -180 -59 -178 -55
rect -152 -59 -150 -56
rect -143 -59 -141 -47
rect -180 -91 -178 -79
rect -152 -92 -150 -79
rect -143 -85 -141 -79
rect -143 -92 -141 -88
rect -180 -105 -178 -101
rect -152 -105 -150 -102
rect -143 -104 -141 -102
rect -142 -108 -141 -104
rect -143 -109 -141 -108
<< polycontact >>
rect -147 -52 -143 -48
rect -178 -90 -174 -86
rect -156 -90 -152 -86
rect -146 -108 -142 -104
<< metal1 >>
rect -192 -50 -173 -47
rect -177 -59 -173 -50
rect -162 -49 -159 -47
rect -162 -52 -147 -49
rect -162 -59 -159 -52
rect -170 -62 -157 -59
rect -185 -95 -182 -79
rect -170 -86 -167 -62
rect -148 -80 -145 -77
rect -174 -89 -167 -86
rect -159 -90 -156 -87
rect -148 -92 -145 -85
rect -186 -97 -182 -95
rect -140 -86 -137 -79
rect -128 -86 -125 -48
rect -140 -88 -125 -86
rect -140 -89 -133 -88
rect -140 -92 -137 -89
rect -128 -89 -125 -88
rect -186 -100 -185 -97
rect -176 -106 -173 -101
rect -192 -109 -173 -106
rect -163 -103 -157 -99
rect -158 -105 -157 -103
rect -158 -108 -146 -105
<< m2contact >>
rect -149 -85 -144 -80
rect -191 -100 -186 -95
rect -163 -108 -158 -103
<< metal2 >>
rect -144 -84 -128 -81
rect -190 -110 -187 -100
rect -163 -110 -160 -108
rect -190 -113 -160 -110
<< m123contact >>
rect -164 -91 -159 -86
rect -133 -93 -128 -88
<< metal3 >>
rect -159 -88 -130 -87
rect -159 -90 -133 -88
<< labels >>
rlabel metal3 -135 -87 -135 -87 1 in2
rlabel m2contact -161 -107 -161 -107 1 in1_inv
rlabel metal1 -170 -89 -167 -87 7 in1
rlabel metal1 -177 -108 -177 -108 1 gnd
rlabel metal1 -186 -49 -186 -49 5 vdd
rlabel metal1 -148 -87 -146 -85 1 s1
<< end >>
