magic
tech scmos
timestamp 1731417668
<< nwell >>
rect 396 149 473 171
rect 513 165 545 184
rect 378 139 473 149
rect 491 159 545 165
rect 378 119 430 139
rect 491 131 543 159
rect 378 117 402 119
rect 481 71 515 123
rect 532 111 566 117
rect 532 85 588 111
rect 563 79 588 85
<< ntransistor >>
rect 551 170 561 172
rect 555 152 565 154
rect 555 142 565 144
rect 389 101 391 111
rect 450 107 452 127
rect 460 107 462 127
rect 407 97 409 107
rect 417 97 419 107
rect 492 49 494 59
rect 502 49 504 59
rect 543 53 545 73
rect 553 53 555 73
rect 574 63 576 73
<< ptransistor >>
rect 519 170 539 172
rect 389 123 391 143
rect 407 125 409 165
rect 417 125 419 165
rect 450 145 452 165
rect 460 145 462 165
rect 497 152 537 154
rect 497 142 537 144
rect 492 77 494 117
rect 502 77 504 117
rect 543 91 545 111
rect 553 91 555 111
rect 574 85 576 105
<< ndiffusion >>
rect 555 173 561 177
rect 551 172 561 173
rect 551 169 561 170
rect 551 165 557 169
rect 555 155 561 159
rect 555 154 565 155
rect 555 150 565 152
rect 559 146 565 150
rect 555 144 565 146
rect 555 141 565 142
rect 555 137 561 141
rect 388 107 389 111
rect 384 101 389 107
rect 391 105 396 111
rect 449 123 450 127
rect 445 107 450 123
rect 452 107 460 127
rect 462 111 467 127
rect 462 107 463 111
rect 391 101 392 105
rect 402 101 407 107
rect 406 97 407 101
rect 409 103 411 107
rect 415 103 417 107
rect 409 97 417 103
rect 419 101 424 107
rect 419 97 420 101
rect 487 53 492 59
rect 491 49 492 53
rect 494 55 496 59
rect 500 55 502 59
rect 494 49 502 55
rect 504 53 509 59
rect 538 57 543 73
rect 542 53 543 57
rect 545 53 553 73
rect 555 69 556 73
rect 555 53 560 69
rect 569 67 574 73
rect 573 63 574 67
rect 576 69 577 73
rect 576 63 581 69
rect 504 49 505 53
<< pdiffusion >>
rect 519 173 535 177
rect 519 172 539 173
rect 519 169 539 170
rect 523 165 539 169
rect 384 127 389 143
rect 388 123 389 127
rect 391 139 392 143
rect 391 123 396 139
rect 402 129 407 165
rect 406 125 407 129
rect 409 125 417 165
rect 419 161 420 165
rect 419 125 424 161
rect 449 161 450 165
rect 445 145 450 161
rect 452 149 460 165
rect 452 145 454 149
rect 458 145 460 149
rect 462 161 463 165
rect 462 145 467 161
rect 497 155 533 159
rect 497 154 537 155
rect 497 144 537 152
rect 497 141 537 142
rect 501 137 537 141
rect 491 113 492 117
rect 487 77 492 113
rect 494 77 502 117
rect 504 81 509 117
rect 542 107 543 111
rect 538 91 543 107
rect 545 95 553 111
rect 545 91 547 95
rect 551 91 553 95
rect 555 107 556 111
rect 555 91 560 107
rect 573 101 574 105
rect 504 77 505 81
rect 569 85 574 101
rect 576 89 581 105
rect 576 85 577 89
<< ndcontact >>
rect 551 173 555 177
rect 557 165 561 169
rect 561 155 565 159
rect 555 146 559 150
rect 561 137 565 141
rect 384 107 388 111
rect 445 123 449 127
rect 463 107 467 111
rect 392 101 396 105
rect 402 97 406 101
rect 411 103 415 107
rect 420 97 424 101
rect 487 49 491 53
rect 496 55 500 59
rect 538 53 542 57
rect 556 69 560 73
rect 569 63 573 67
rect 577 69 581 73
rect 505 49 509 53
<< pdcontact >>
rect 535 173 539 177
rect 519 165 523 169
rect 384 123 388 127
rect 392 139 396 143
rect 402 125 406 129
rect 420 161 424 165
rect 445 161 449 165
rect 454 145 458 149
rect 463 161 467 165
rect 533 155 537 159
rect 497 137 501 141
rect 487 113 491 117
rect 538 107 542 111
rect 547 91 551 95
rect 556 107 560 111
rect 569 101 573 105
rect 505 77 509 81
rect 577 85 581 89
<< polysilicon >>
rect 516 170 519 172
rect 539 170 551 172
rect 561 170 564 172
rect 407 165 409 168
rect 417 165 419 168
rect 450 165 452 169
rect 460 165 462 169
rect 389 143 391 146
rect 494 152 497 154
rect 537 152 555 154
rect 565 152 568 154
rect 450 127 452 145
rect 460 127 462 145
rect 494 142 497 144
rect 537 142 555 144
rect 565 142 568 144
rect 389 111 391 123
rect 407 107 409 125
rect 417 107 419 125
rect 492 117 494 120
rect 502 117 504 120
rect 389 98 391 101
rect 450 103 452 107
rect 460 103 462 107
rect 407 94 409 97
rect 417 94 419 97
rect 543 111 545 115
rect 553 111 555 115
rect 574 105 576 109
rect 492 59 494 77
rect 502 59 504 77
rect 543 73 545 91
rect 553 73 555 91
rect 574 73 576 85
rect 574 59 576 63
rect 543 49 545 53
rect 553 49 555 53
rect 492 46 494 49
rect 502 46 504 49
<< polycontact >>
rect 546 166 550 170
rect 452 128 456 132
rect 544 148 548 152
rect 462 134 466 138
rect 550 138 554 142
rect 391 112 395 116
rect 409 114 413 118
rect 419 108 423 112
rect 539 80 543 84
rect 488 60 492 64
rect 498 66 502 70
rect 549 74 553 78
rect 570 74 574 78
<< metal1 >>
rect 509 181 549 184
rect 393 172 468 175
rect 509 175 512 181
rect 546 177 549 181
rect 481 172 512 175
rect 539 174 551 177
rect 393 143 396 172
rect 421 165 424 172
rect 445 165 449 172
rect 464 165 467 172
rect 454 144 457 145
rect 445 141 457 144
rect 445 132 448 141
rect 481 138 484 172
rect 466 135 484 138
rect 492 165 519 168
rect 487 140 490 163
rect 546 159 549 166
rect 561 165 572 168
rect 569 159 572 165
rect 537 156 554 159
rect 551 150 554 156
rect 565 156 572 159
rect 487 137 497 140
rect 427 129 448 132
rect 384 116 387 123
rect 402 116 405 125
rect 427 118 430 129
rect 445 127 448 129
rect 456 128 473 131
rect 487 127 490 137
rect 544 131 547 148
rect 551 147 555 150
rect 569 141 572 156
rect 550 131 553 138
rect 565 137 569 140
rect 487 124 535 127
rect 377 113 387 116
rect 384 111 387 113
rect 395 113 405 116
rect 413 115 430 118
rect 487 117 490 124
rect 532 121 535 124
rect 532 118 572 121
rect 402 111 405 113
rect 402 108 414 111
rect 423 109 427 112
rect 411 107 414 108
rect 538 111 541 118
rect 556 111 560 118
rect 464 102 467 107
rect 569 105 572 118
rect 393 93 396 101
rect 402 93 405 97
rect 421 93 424 97
rect 428 99 476 102
rect 428 93 431 99
rect 393 90 431 93
rect 473 45 476 99
rect 548 90 551 91
rect 548 87 560 90
rect 512 81 539 84
rect 485 67 498 70
rect 506 68 509 77
rect 512 68 515 81
rect 557 78 560 87
rect 578 78 581 85
rect 532 74 549 77
rect 557 75 570 78
rect 557 73 560 75
rect 578 75 584 78
rect 578 73 581 75
rect 506 65 515 68
rect 480 61 488 64
rect 506 63 509 65
rect 497 60 509 63
rect 497 59 500 60
rect 487 45 490 49
rect 506 45 509 49
rect 538 48 541 53
rect 569 49 572 63
rect 532 45 568 48
rect 473 42 536 45
<< m2contact >>
rect 468 172 473 177
rect 487 163 492 168
rect 542 126 547 131
rect 480 67 485 72
rect 584 73 589 78
rect 479 56 484 61
<< metal2 >>
rect 473 173 490 176
rect 487 168 490 173
rect 480 127 542 130
rect 480 72 483 127
rect 529 112 588 115
rect 585 78 588 112
<< m3contact >>
rect 524 111 529 116
<< m123contact >>
rect 569 136 574 141
rect 427 107 432 112
rect 568 44 573 49
<< metal3 >>
rect 523 116 530 117
rect 523 115 524 116
rect 431 112 524 115
rect 432 109 434 112
rect 523 111 524 112
rect 529 111 530 116
rect 523 110 530 111
rect 570 49 573 136
<< labels >>
rlabel metal1 488 125 488 126 5 vdd
rlabel metal1 498 44 498 44 1 gnd
rlabel metal1 544 119 544 119 5 vdd
rlabel metal1 553 46 553 46 1 gnd
rlabel metal1 570 148 570 148 7 gnd
rlabel metal1 488 138 489 138 3 vdd
rlabel metal1 461 173 461 173 5 vdd
rlabel metal1 452 100 452 100 1 gnd
rlabel metal1 423 173 423 174 5 vdd
rlabel metal1 413 92 413 92 1 gnd
rlabel metal1 384 114 386 116 1 c3
rlabel metal1 439 129 445 132 1 temp108
rlabel metal1 579 76 581 78 1 temp106
rlabel metal1 533 75 537 76 1 c1
rlabel metal1 510 65 514 67 1 temp105
rlabel metal1 550 132 553 135 1 g1_inv
rlabel metal1 483 67 487 69 1 p2_inv
rlabel metal1 545 174 548 177 1 temp107
rlabel metal1 481 61 486 63 1 p1_inv
rlabel metal1 468 128 470 130 1 g2_inv
<< end >>
