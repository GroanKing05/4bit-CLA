magic
tech scmos
timestamp 1731426146
<< nwell >>
rect -118 70 -84 90
rect -118 68 -50 70
rect -137 64 -50 68
rect -137 38 -29 64
rect -137 36 -112 38
rect -53 32 -29 38
rect -18 58 16 80
rect -18 28 35 58
rect 10 26 35 28
rect 41 26 75 58
rect -37 -46 15 -12
<< ntransistor >>
rect -125 20 -123 30
rect -107 16 -105 26
rect -97 16 -95 26
rect -73 6 -71 26
rect -63 6 -61 26
rect -42 16 -40 26
rect -7 6 -5 16
rect 3 6 5 16
rect 21 10 23 20
rect 52 -6 54 14
rect 62 -6 64 14
rect 27 -25 37 -23
rect 27 -35 37 -33
<< ptransistor >>
rect -125 42 -123 62
rect -107 44 -105 84
rect -97 44 -95 84
rect -73 44 -71 64
rect -63 44 -61 64
rect -42 38 -40 58
rect -7 34 -5 74
rect 3 34 5 74
rect 21 32 23 52
rect 52 32 54 52
rect 62 32 64 52
rect -31 -25 9 -23
rect -31 -35 9 -33
<< ndiffusion >>
rect -126 26 -125 30
rect -130 20 -125 26
rect -123 24 -118 30
rect -123 20 -122 24
rect -112 20 -107 26
rect -108 16 -107 20
rect -105 22 -103 26
rect -99 22 -97 26
rect -105 16 -97 22
rect -95 20 -90 26
rect -95 16 -94 20
rect -78 10 -73 26
rect -74 6 -73 10
rect -71 6 -63 26
rect -61 22 -60 26
rect -61 6 -56 22
rect -47 20 -42 26
rect -43 16 -42 20
rect -40 22 -39 26
rect -40 16 -35 22
rect -12 10 -7 16
rect -8 6 -7 10
rect -5 12 -3 16
rect 1 12 3 16
rect -5 6 3 12
rect 5 10 10 16
rect 16 14 21 20
rect 20 10 21 14
rect 23 16 24 20
rect 23 10 28 16
rect 5 6 6 10
rect 47 -2 52 14
rect 51 -6 52 -2
rect 54 -6 62 14
rect 64 10 65 14
rect 64 -6 69 10
rect 27 -22 33 -18
rect 27 -23 37 -22
rect 27 -27 37 -25
rect 31 -31 37 -27
rect 27 -33 37 -31
rect 27 -36 37 -35
rect 27 -40 33 -36
<< pdiffusion >>
rect -130 46 -125 62
rect -126 42 -125 46
rect -123 58 -122 62
rect -123 42 -118 58
rect -112 48 -107 84
rect -108 44 -107 48
rect -105 44 -97 84
rect -95 80 -94 84
rect -95 44 -90 80
rect -8 70 -7 74
rect -74 60 -73 64
rect -78 44 -73 60
rect -71 48 -63 64
rect -71 44 -69 48
rect -65 44 -63 48
rect -61 60 -60 64
rect -61 44 -56 60
rect -43 54 -42 58
rect -47 38 -42 54
rect -40 42 -35 58
rect -40 38 -39 42
rect -12 34 -7 70
rect -5 34 3 74
rect 5 38 10 74
rect 5 34 6 38
rect 20 48 21 52
rect 16 32 21 48
rect 23 36 28 52
rect 23 32 24 36
rect 51 48 52 52
rect 47 32 52 48
rect 54 36 62 52
rect 54 32 56 36
rect 60 32 62 36
rect 64 48 65 52
rect 64 32 69 48
rect -27 -22 9 -18
rect -31 -23 9 -22
rect -31 -33 9 -25
rect -31 -36 9 -35
rect -31 -40 5 -36
<< ndcontact >>
rect -130 26 -126 30
rect -122 20 -118 24
rect -112 16 -108 20
rect -103 22 -99 26
rect -94 16 -90 20
rect -78 6 -74 10
rect -60 22 -56 26
rect -47 16 -43 20
rect -39 22 -35 26
rect -12 6 -8 10
rect -3 12 1 16
rect 16 10 20 14
rect 24 16 28 20
rect 6 6 10 10
rect 47 -6 51 -2
rect 65 10 69 14
rect 33 -22 37 -18
rect 27 -31 31 -27
rect 33 -40 37 -36
<< pdcontact >>
rect -130 42 -126 46
rect -122 58 -118 62
rect -112 44 -108 48
rect -94 80 -90 84
rect -12 70 -8 74
rect -78 60 -74 64
rect -69 44 -65 48
rect -60 60 -56 64
rect -47 54 -43 58
rect -39 38 -35 42
rect 6 34 10 38
rect 16 48 20 52
rect 24 32 28 36
rect 47 48 51 52
rect 56 32 60 36
rect 65 48 69 52
rect -31 -22 -27 -18
rect 5 -40 9 -36
<< polysilicon >>
rect -107 84 -105 87
rect -97 84 -95 87
rect -125 62 -123 65
rect -7 74 -5 77
rect 3 74 5 77
rect -73 64 -71 68
rect -63 64 -61 68
rect -42 58 -40 62
rect -125 30 -123 42
rect -107 26 -105 44
rect -97 26 -95 44
rect -73 26 -71 44
rect -63 26 -61 44
rect -42 26 -40 38
rect 21 52 23 55
rect 52 52 54 56
rect 62 52 64 56
rect -125 17 -123 20
rect -107 13 -105 16
rect -97 13 -95 16
rect -7 16 -5 34
rect 3 16 5 34
rect 21 20 23 32
rect -42 12 -40 16
rect 52 14 54 32
rect 62 14 64 32
rect 21 7 23 10
rect -73 2 -71 6
rect -63 2 -61 6
rect -7 3 -5 6
rect 3 3 5 6
rect 52 -10 54 -6
rect 62 -10 64 -6
rect -34 -25 -31 -23
rect 9 -25 27 -23
rect 37 -25 40 -23
rect -34 -35 -31 -33
rect 9 -35 27 -33
rect 37 -35 40 -33
<< polycontact >>
rect -123 31 -119 35
rect -105 33 -101 37
rect -77 34 -73 38
rect -95 27 -91 31
rect -67 27 -63 31
rect -46 27 -42 31
rect -11 17 -7 21
rect -1 23 3 27
rect 17 21 21 25
rect 48 21 52 25
rect 58 15 62 19
rect 22 -23 26 -19
rect 16 -33 20 -29
<< metal1 >>
rect -121 91 -80 94
rect -121 72 -118 91
rect -93 84 -90 91
rect -132 69 -118 72
rect -83 74 -80 91
rect -47 81 19 84
rect -47 74 -44 81
rect -83 71 -44 74
rect -121 62 -118 69
rect -78 64 -75 71
rect -60 64 -56 71
rect -47 58 -44 71
rect -12 74 -9 81
rect 16 62 19 81
rect 16 59 75 62
rect 16 52 19 59
rect 47 52 50 59
rect 65 52 69 59
rect -130 35 -127 42
rect -112 35 -109 44
rect -68 43 -65 44
rect -68 40 -56 43
rect -137 32 -127 35
rect -130 30 -127 32
rect -119 32 -109 35
rect -101 34 -77 37
rect -112 30 -109 32
rect -59 31 -56 40
rect -38 31 -35 38
rect -112 27 -100 30
rect -91 28 -67 31
rect -59 28 -46 31
rect -103 26 -100 27
rect -59 26 -56 28
rect -38 26 -31 31
rect -35 22 -31 26
rect -14 24 -1 27
rect 7 25 10 34
rect 25 25 28 32
rect 57 31 60 32
rect 57 28 69 31
rect -121 12 -118 20
rect -112 12 -109 16
rect -93 12 -90 16
rect -121 9 -82 12
rect -85 1 -82 9
rect -78 1 -75 6
rect -47 2 -44 16
rect -34 13 -31 22
rect 7 22 17 25
rect -19 19 -11 20
rect -14 17 -11 19
rect 7 20 10 22
rect 25 22 48 25
rect 25 20 28 22
rect -2 17 10 20
rect -2 16 1 17
rect 66 19 69 28
rect -33 8 -31 13
rect 41 15 58 18
rect 66 16 79 19
rect 66 14 69 16
rect -12 2 -9 6
rect 7 2 10 6
rect 16 2 19 10
rect -47 1 44 2
rect -85 -1 44 1
rect -85 -2 -44 -1
rect -41 -18 -38 -16
rect -41 -21 -31 -18
rect -41 -46 -38 -21
rect 16 -29 19 -4
rect 41 -11 44 -1
rect 76 -4 79 16
rect 47 -11 50 -6
rect 41 -14 72 -11
rect 22 -19 25 -14
rect 41 -18 44 -14
rect 37 -21 44 -18
rect 23 -31 27 -28
rect 23 -37 26 -31
rect 9 -40 26 -37
rect 41 -37 44 -21
rect 37 -40 44 -37
rect 18 -46 21 -40
<< m2contact >>
rect -19 23 -14 28
rect -19 14 -14 19
rect -38 8 -33 13
rect 11 -9 16 -4
rect 22 -14 27 -9
rect 76 -9 81 -4
<< metal2 >>
rect -37 -3 -34 8
rect -37 -4 16 -3
rect -37 -6 11 -4
rect 22 -8 76 -5
rect 22 -9 27 -8
<< m123contact >>
rect -137 69 -132 74
rect -43 -16 -38 -11
<< metal3 >>
rect -136 16 -133 69
rect -136 13 -122 16
rect -125 7 -122 13
rect -125 4 -86 7
rect -89 -4 -86 4
rect -89 -7 -39 -4
rect -42 -11 -39 -7
<< labels >>
rlabel metal1 -72 72 -72 72 5 vdd
rlabel metal1 -63 -1 -63 -1 1 gnd
rlabel metal1 -36 29 -36 31 1 temp110
rlabel metal1 -101 11 -101 11 1 gnd
rlabel metal1 -91 92 -91 93 5 vdd
rlabel metal1 -84 29 -84 29 1 temp109
rlabel metal1 -90 34 -78 37 1 temp104
rlabel metal1 -130 33 -130 33 1 temp110
rlabel metal1 -11 82 -11 83 5 vdd
rlabel metal1 -1 1 -1 1 1 gnd
rlabel metal1 26 23 28 25 1 temp111
rlabel m2contact -17 24 -14 26 1 g2_inv
rlabel m2contact -15 17 -15 17 1 p3_inv
rlabel metal1 53 60 53 60 5 vdd
rlabel metal1 62 -13 62 -13 1 gnd
rlabel metal1 43 15 45 18 1 g3_inv
rlabel metal1 69 16 75 19 7 temp112
rlabel metal1 -40 -19 -39 -19 3 vdd
rlabel metal1 42 -29 42 -29 7 gnd
rlabel metal1 19 -45 21 -42 1 g4_inv
<< end >>
