magic
tech scmos
timestamp 1731623447
<< nwell >>
rect -629 -352 -597 -185
rect -529 -314 -497 -147
rect -327 -194 -295 -27
rect -124 -106 -92 61
rect -196 -163 -119 -141
rect -79 -147 -47 -128
rect -214 -173 -119 -163
rect -101 -153 -47 -147
rect -214 -193 -162 -173
rect -101 -181 -49 -153
rect -214 -195 -190 -193
rect -382 -228 -350 -209
rect -382 -234 -328 -228
rect -380 -262 -328 -234
rect -310 -244 -233 -222
rect -111 -241 -77 -189
rect -60 -201 -26 -195
rect -60 -227 -4 -201
rect -29 -233 -4 -227
rect 19 -237 51 -70
rect -310 -254 -215 -244
rect -403 -282 -369 -276
rect -425 -308 -369 -282
rect -425 -314 -400 -308
rect -352 -322 -318 -270
rect -267 -274 -215 -254
rect -239 -276 -215 -274
rect 14 -275 48 -255
rect 14 -277 82 -275
rect -5 -281 82 -277
rect -5 -307 103 -281
rect -5 -309 20 -307
rect 79 -313 103 -307
rect 114 -287 148 -265
rect 114 -317 167 -287
rect -545 -363 -487 -341
rect -285 -350 -224 -318
rect 142 -319 167 -317
rect 173 -319 207 -287
rect -145 -329 -111 -324
rect -182 -335 -111 -329
rect -204 -361 -111 -335
rect -545 -373 -438 -363
rect -204 -367 -179 -361
rect -616 -414 -555 -382
rect -521 -393 -438 -373
rect -493 -395 -438 -393
rect -422 -402 -361 -370
rect -145 -376 -111 -361
rect -90 -392 -29 -360
rect 95 -391 147 -357
rect 43 -432 111 -400
rect -261 -467 -200 -466
rect -109 -467 -48 -466
rect -570 -470 -509 -469
rect -410 -470 -349 -469
rect -570 -481 -472 -470
rect -410 -481 -312 -470
rect -261 -478 -163 -467
rect -109 -478 -11 -467
rect -570 -501 -438 -481
rect -410 -501 -278 -481
rect -261 -498 -129 -478
rect -109 -498 23 -478
rect -506 -513 -438 -501
rect -346 -513 -278 -501
rect -197 -510 -129 -498
rect -45 -510 23 -498
rect -506 -522 -472 -513
rect -346 -522 -312 -513
rect -197 -519 -163 -510
rect -45 -519 -11 -510
rect -614 -680 -582 -538
rect -535 -681 -503 -539
rect -453 -678 -421 -536
rect -369 -679 -337 -537
rect -287 -678 -255 -536
rect -201 -678 -169 -536
rect -116 -679 -84 -537
rect -33 -679 -1 -537
rect 51 -679 83 -537
<< ntransistor >>
rect -86 47 -76 49
rect -82 23 -72 25
rect -86 7 -66 9
rect -86 -2 -66 0
rect -86 -18 -66 -16
rect -86 -27 -66 -25
rect -289 -41 -279 -39
rect -82 -45 -72 -43
rect -285 -65 -275 -63
rect -86 -71 -66 -69
rect -289 -81 -269 -79
rect 57 -84 67 -82
rect -289 -90 -269 -88
rect -86 -95 -66 -93
rect -289 -106 -269 -104
rect 61 -108 71 -106
rect -289 -115 -269 -113
rect 57 -124 77 -122
rect -285 -133 -275 -131
rect 57 -133 77 -131
rect -41 -142 -31 -140
rect -289 -159 -269 -157
rect -491 -161 -481 -159
rect -289 -183 -269 -181
rect -487 -185 -477 -183
rect 57 -149 77 -147
rect 57 -158 77 -156
rect -37 -160 -27 -158
rect -37 -170 -27 -168
rect 61 -176 71 -174
rect -591 -199 -581 -197
rect -491 -201 -471 -199
rect -491 -210 -471 -208
rect -203 -211 -201 -201
rect -142 -205 -140 -185
rect -132 -205 -130 -185
rect -185 -215 -183 -205
rect -175 -215 -173 -205
rect -587 -223 -577 -221
rect -398 -223 -388 -221
rect -491 -226 -471 -224
rect -491 -235 -471 -233
rect -591 -239 -571 -237
rect -402 -241 -392 -239
rect -591 -248 -571 -246
rect -402 -251 -392 -249
rect -487 -253 -477 -251
rect -591 -264 -571 -262
rect -591 -273 -571 -271
rect -491 -279 -471 -277
rect -587 -291 -577 -289
rect -491 -303 -471 -301
rect -591 -317 -571 -315
rect -299 -286 -297 -266
rect -289 -286 -287 -266
rect 57 -202 77 -200
rect 57 -226 77 -224
rect -100 -263 -98 -253
rect -90 -263 -88 -253
rect -49 -259 -47 -239
rect -39 -259 -37 -239
rect -18 -249 -16 -239
rect -256 -296 -254 -286
rect -246 -296 -244 -286
rect -228 -292 -226 -282
rect -413 -330 -411 -320
rect -591 -341 -571 -339
rect -392 -340 -390 -320
rect -382 -340 -380 -320
rect -341 -344 -339 -334
rect -331 -344 -329 -334
rect 7 -325 9 -315
rect 25 -329 27 -319
rect 35 -329 37 -319
rect -534 -389 -532 -379
rect -274 -367 -272 -357
rect -265 -367 -263 -357
rect -237 -366 -235 -356
rect 59 -339 61 -319
rect 69 -339 71 -319
rect 90 -329 92 -319
rect 125 -339 127 -329
rect 135 -339 137 -329
rect 153 -335 155 -325
rect 184 -351 186 -331
rect 194 -351 196 -331
rect -510 -415 -508 -405
rect -500 -415 -498 -405
rect -482 -411 -480 -401
rect -192 -383 -190 -373
rect -171 -393 -169 -373
rect -161 -393 -159 -373
rect 159 -370 169 -368
rect 159 -380 169 -378
rect -605 -431 -603 -421
rect -596 -431 -594 -421
rect -568 -430 -566 -420
rect -461 -427 -459 -407
rect -451 -427 -449 -407
rect -134 -398 -132 -388
rect -124 -398 -122 -388
rect -79 -408 -77 -398
rect -411 -419 -409 -409
rect -402 -419 -400 -409
rect -374 -418 -372 -408
rect -51 -409 -49 -399
rect -42 -409 -40 -399
rect -559 -462 -557 -452
rect -550 -462 -548 -452
rect -522 -463 -520 -453
rect -495 -458 -493 -448
rect -485 -458 -483 -448
rect -461 -469 -459 -449
rect -451 -469 -449 -449
rect -399 -462 -397 -452
rect -390 -462 -388 -452
rect -362 -463 -360 -453
rect -335 -458 -333 -448
rect -325 -458 -323 -448
rect -301 -469 -299 -449
rect -291 -469 -289 -449
rect -250 -459 -248 -449
rect -241 -459 -239 -449
rect -213 -460 -211 -450
rect -186 -455 -184 -445
rect -176 -455 -174 -445
rect -152 -466 -150 -446
rect -142 -466 -140 -446
rect -98 -459 -96 -449
rect -89 -459 -87 -449
rect -61 -460 -59 -450
rect -34 -455 -32 -445
rect -24 -455 -22 -445
rect 0 -466 2 -446
rect 10 -466 12 -446
rect 54 -464 56 -444
rect 64 -464 66 -444
rect 88 -464 90 -444
rect 98 -464 100 -444
rect -572 -551 -562 -549
rect -411 -549 -401 -547
rect -493 -552 -483 -550
rect -327 -550 -317 -548
rect -245 -549 -235 -547
rect -159 -549 -149 -547
rect -74 -550 -64 -548
rect 9 -550 19 -548
rect 93 -550 103 -548
rect -415 -565 -395 -563
rect -576 -567 -556 -565
rect -497 -568 -477 -566
rect -576 -576 -556 -574
rect -331 -566 -311 -564
rect -249 -565 -229 -563
rect -163 -565 -143 -563
rect -415 -574 -395 -572
rect -78 -566 -58 -564
rect 5 -566 25 -564
rect 89 -566 109 -564
rect -497 -577 -477 -575
rect -331 -575 -311 -573
rect -249 -574 -229 -572
rect -163 -574 -143 -572
rect -78 -575 -58 -573
rect 5 -575 25 -573
rect 89 -575 109 -573
rect -415 -590 -395 -588
rect -576 -592 -556 -590
rect -497 -593 -477 -591
rect -576 -601 -556 -599
rect -331 -591 -311 -589
rect -249 -590 -229 -588
rect -163 -590 -143 -588
rect -415 -599 -395 -597
rect -78 -591 -58 -589
rect 5 -591 25 -589
rect 89 -591 109 -589
rect -497 -602 -477 -600
rect -331 -600 -311 -598
rect -249 -599 -229 -597
rect -163 -599 -143 -597
rect -78 -600 -58 -598
rect 5 -600 25 -598
rect 89 -600 109 -598
rect -572 -619 -562 -617
rect -411 -617 -401 -615
rect -493 -620 -483 -618
rect -327 -618 -317 -616
rect -245 -617 -235 -615
rect -159 -617 -149 -615
rect -74 -618 -64 -616
rect 9 -618 19 -616
rect 93 -618 103 -616
rect -576 -645 -556 -643
rect -415 -643 -395 -641
rect -497 -646 -477 -644
rect -331 -644 -311 -642
rect -249 -643 -229 -641
rect -163 -643 -143 -641
rect -78 -644 -58 -642
rect 5 -644 25 -642
rect 89 -644 109 -642
rect -576 -669 -556 -667
rect -415 -667 -395 -665
rect -497 -670 -477 -668
rect -331 -668 -311 -666
rect -249 -667 -229 -665
rect -163 -667 -143 -665
rect -78 -668 -58 -666
rect 5 -668 25 -666
rect 89 -668 109 -666
<< ptransistor >>
rect -118 47 -98 49
rect -118 23 -98 25
rect -118 -2 -98 0
rect -118 -27 -98 -25
rect -321 -41 -301 -39
rect -118 -45 -98 -43
rect -118 -63 -98 -61
rect -321 -65 -301 -63
rect -118 -71 -98 -69
rect 25 -84 45 -82
rect -118 -87 -98 -85
rect -321 -90 -301 -88
rect -118 -95 -98 -93
rect 25 -108 45 -106
rect -321 -115 -301 -113
rect -321 -133 -301 -131
rect 25 -133 45 -131
rect -73 -142 -53 -140
rect -321 -151 -301 -149
rect -321 -159 -301 -157
rect -523 -161 -503 -159
rect -321 -175 -301 -173
rect -321 -183 -301 -181
rect -523 -185 -503 -183
rect -203 -189 -201 -169
rect -185 -187 -183 -147
rect -175 -187 -173 -147
rect -142 -167 -140 -147
rect -132 -167 -130 -147
rect 25 -158 45 -156
rect -95 -160 -55 -158
rect -95 -170 -55 -168
rect 25 -176 45 -174
rect -623 -199 -603 -197
rect -523 -210 -503 -208
rect 25 -194 45 -192
rect -623 -223 -603 -221
rect -376 -223 -356 -221
rect -523 -235 -503 -233
rect -374 -241 -334 -239
rect -623 -248 -603 -246
rect -299 -248 -297 -228
rect -289 -248 -287 -228
rect -374 -251 -334 -249
rect -523 -253 -503 -251
rect -523 -271 -503 -269
rect -623 -273 -603 -271
rect -523 -279 -503 -277
rect -623 -291 -603 -289
rect -523 -295 -503 -293
rect -523 -303 -503 -301
rect -623 -309 -603 -307
rect -413 -308 -411 -288
rect -392 -302 -390 -282
rect -382 -302 -380 -282
rect -623 -317 -603 -315
rect -341 -316 -339 -276
rect -331 -316 -329 -276
rect -256 -268 -254 -228
rect -246 -268 -244 -228
rect -100 -235 -98 -195
rect -90 -235 -88 -195
rect -49 -221 -47 -201
rect -39 -221 -37 -201
rect 25 -202 45 -200
rect -228 -270 -226 -250
rect -18 -227 -16 -207
rect 25 -218 45 -216
rect 25 -226 45 -224
rect 7 -303 9 -283
rect 25 -301 27 -261
rect 35 -301 37 -261
rect 59 -301 61 -281
rect 69 -301 71 -281
rect -623 -333 -603 -331
rect -623 -341 -603 -339
rect -274 -344 -272 -324
rect -265 -344 -263 -324
rect -237 -344 -235 -324
rect 90 -307 92 -287
rect 125 -311 127 -271
rect 135 -311 137 -271
rect -534 -367 -532 -347
rect -605 -408 -603 -388
rect -596 -408 -594 -388
rect -568 -408 -566 -388
rect -510 -387 -508 -347
rect -500 -387 -498 -347
rect -482 -389 -480 -369
rect -461 -389 -459 -369
rect -451 -389 -449 -369
rect -192 -361 -190 -341
rect -171 -355 -169 -335
rect -161 -355 -159 -335
rect -134 -370 -132 -330
rect -124 -370 -122 -330
rect 153 -313 155 -293
rect 184 -313 186 -293
rect 194 -313 196 -293
rect -411 -396 -409 -376
rect -402 -396 -400 -376
rect -374 -396 -372 -376
rect -79 -386 -77 -366
rect -51 -386 -49 -366
rect -42 -386 -40 -366
rect 101 -370 141 -368
rect 101 -380 141 -378
rect 54 -426 56 -406
rect 64 -426 66 -406
rect 88 -426 90 -406
rect 98 -426 100 -406
rect -559 -495 -557 -475
rect -550 -495 -548 -475
rect -522 -495 -520 -475
rect -495 -516 -493 -476
rect -485 -516 -483 -476
rect -461 -507 -459 -487
rect -451 -507 -449 -487
rect -399 -495 -397 -475
rect -390 -495 -388 -475
rect -362 -495 -360 -475
rect -335 -516 -333 -476
rect -325 -516 -323 -476
rect -301 -507 -299 -487
rect -291 -507 -289 -487
rect -250 -492 -248 -472
rect -241 -492 -239 -472
rect -213 -492 -211 -472
rect -186 -513 -184 -473
rect -176 -513 -174 -473
rect -152 -504 -150 -484
rect -142 -504 -140 -484
rect -98 -492 -96 -472
rect -89 -492 -87 -472
rect -61 -492 -59 -472
rect -34 -513 -32 -473
rect -24 -513 -22 -473
rect 0 -504 2 -484
rect 10 -504 12 -484
rect -608 -551 -588 -549
rect -447 -549 -427 -547
rect -529 -552 -509 -550
rect -363 -550 -343 -548
rect -281 -549 -261 -547
rect -195 -549 -175 -547
rect -110 -550 -90 -548
rect -27 -550 -7 -548
rect 57 -550 77 -548
rect -608 -576 -588 -574
rect -447 -574 -427 -572
rect -529 -577 -509 -575
rect -363 -575 -343 -573
rect -281 -574 -261 -572
rect -195 -574 -175 -572
rect -110 -575 -90 -573
rect -27 -575 -7 -573
rect 57 -575 77 -573
rect -608 -601 -588 -599
rect -447 -599 -427 -597
rect -529 -602 -509 -600
rect -363 -600 -343 -598
rect -281 -599 -261 -597
rect -195 -599 -175 -597
rect -110 -600 -90 -598
rect -27 -600 -7 -598
rect 57 -600 77 -598
rect -608 -619 -588 -617
rect -447 -617 -427 -615
rect -529 -620 -509 -618
rect -363 -618 -343 -616
rect -281 -617 -261 -615
rect -195 -617 -175 -615
rect -110 -618 -90 -616
rect -27 -618 -7 -616
rect 57 -618 77 -616
rect -447 -635 -427 -633
rect -608 -637 -588 -635
rect -529 -638 -509 -636
rect -608 -645 -588 -643
rect -363 -636 -343 -634
rect -281 -635 -261 -633
rect -195 -635 -175 -633
rect -447 -643 -427 -641
rect -110 -636 -90 -634
rect -27 -636 -7 -634
rect 57 -636 77 -634
rect -529 -646 -509 -644
rect -363 -644 -343 -642
rect -281 -643 -261 -641
rect -195 -643 -175 -641
rect -110 -644 -90 -642
rect -27 -644 -7 -642
rect 57 -644 77 -642
rect -447 -659 -427 -657
rect -608 -661 -588 -659
rect -529 -662 -509 -660
rect -608 -669 -588 -667
rect -363 -660 -343 -658
rect -281 -659 -261 -657
rect -447 -667 -427 -665
rect -195 -659 -175 -657
rect -110 -660 -90 -658
rect -529 -670 -509 -668
rect -363 -668 -343 -666
rect -281 -667 -261 -665
rect -195 -667 -175 -665
rect -27 -660 -7 -658
rect 57 -660 77 -658
rect -110 -668 -90 -666
rect -27 -668 -7 -666
rect 57 -668 77 -666
<< ndiffusion >>
rect -82 50 -76 54
rect -86 49 -76 50
rect -86 46 -76 47
rect -86 42 -80 46
rect -78 26 -72 30
rect -82 25 -72 26
rect -82 22 -72 23
rect -82 18 -76 22
rect -82 10 -66 14
rect -86 9 -66 10
rect -86 0 -66 7
rect -86 -3 -66 -2
rect -86 -7 -70 -3
rect -82 -15 -66 -11
rect -86 -16 -66 -15
rect -86 -25 -66 -18
rect -86 -28 -66 -27
rect -86 -32 -70 -28
rect -285 -38 -279 -34
rect -289 -39 -279 -38
rect -289 -42 -279 -41
rect -289 -46 -283 -42
rect -78 -42 -72 -38
rect -82 -43 -72 -42
rect -82 -46 -72 -45
rect -82 -50 -76 -46
rect -281 -62 -275 -58
rect -285 -63 -275 -62
rect -285 -66 -275 -65
rect -285 -70 -279 -66
rect -82 -68 -66 -64
rect -86 -69 -66 -68
rect -285 -78 -269 -74
rect -86 -72 -66 -71
rect -86 -76 -70 -72
rect -289 -79 -269 -78
rect -289 -88 -269 -81
rect 61 -81 67 -77
rect 57 -82 67 -81
rect -289 -91 -269 -90
rect -289 -95 -273 -91
rect -82 -92 -66 -88
rect 57 -85 67 -84
rect 57 -89 63 -85
rect -86 -93 -66 -92
rect -285 -103 -269 -99
rect -86 -96 -66 -95
rect -86 -100 -70 -96
rect -289 -104 -269 -103
rect 65 -105 71 -101
rect 61 -106 71 -105
rect -289 -113 -269 -106
rect 61 -109 71 -108
rect 61 -113 67 -109
rect -289 -116 -269 -115
rect -289 -120 -273 -116
rect 61 -121 77 -117
rect 57 -122 77 -121
rect -281 -130 -275 -126
rect -285 -131 -275 -130
rect 57 -131 77 -124
rect -285 -134 -275 -133
rect -285 -138 -279 -134
rect -37 -139 -31 -135
rect 57 -134 77 -133
rect 57 -138 73 -134
rect -41 -140 -31 -139
rect -41 -143 -31 -142
rect -41 -147 -35 -143
rect 61 -146 77 -142
rect 57 -147 77 -146
rect -487 -158 -481 -154
rect -285 -156 -269 -152
rect -289 -157 -269 -156
rect -491 -159 -481 -158
rect -491 -162 -481 -161
rect -491 -166 -485 -162
rect -289 -160 -269 -159
rect -289 -164 -273 -160
rect -483 -182 -477 -178
rect -285 -180 -269 -176
rect -289 -181 -269 -180
rect -487 -183 -477 -182
rect -487 -186 -477 -185
rect -487 -190 -481 -186
rect -289 -184 -269 -183
rect -289 -188 -273 -184
rect -37 -157 -31 -153
rect 57 -156 77 -149
rect -37 -158 -27 -157
rect -37 -162 -27 -160
rect -33 -166 -27 -162
rect 57 -159 77 -158
rect 57 -163 73 -159
rect -37 -168 -27 -166
rect -37 -171 -27 -170
rect -37 -175 -31 -171
rect 65 -173 71 -169
rect 61 -174 71 -173
rect 61 -177 71 -176
rect 61 -181 67 -177
rect -587 -196 -581 -192
rect -591 -197 -581 -196
rect -487 -198 -471 -194
rect -491 -199 -471 -198
rect -591 -200 -581 -199
rect -591 -204 -585 -200
rect -491 -208 -471 -201
rect -204 -205 -203 -201
rect -491 -211 -471 -210
rect -208 -211 -203 -205
rect -201 -207 -196 -201
rect -143 -189 -142 -185
rect -147 -205 -142 -189
rect -140 -205 -132 -185
rect -130 -201 -125 -185
rect -130 -205 -129 -201
rect -201 -211 -200 -207
rect -190 -211 -185 -205
rect -491 -215 -475 -211
rect -186 -215 -185 -211
rect -183 -209 -181 -205
rect -177 -209 -175 -205
rect -183 -215 -175 -209
rect -173 -211 -168 -205
rect -173 -215 -172 -211
rect -583 -220 -577 -216
rect -587 -221 -577 -220
rect -487 -223 -471 -219
rect -398 -220 -392 -216
rect -398 -221 -388 -220
rect -587 -224 -577 -223
rect -491 -224 -471 -223
rect -398 -224 -388 -223
rect -587 -228 -581 -224
rect -587 -236 -571 -232
rect -491 -233 -471 -226
rect -394 -228 -388 -224
rect -591 -237 -571 -236
rect -591 -246 -571 -239
rect -491 -236 -471 -235
rect -491 -240 -475 -236
rect -398 -238 -392 -234
rect -402 -239 -392 -238
rect -402 -243 -392 -241
rect -591 -249 -571 -248
rect -591 -253 -575 -249
rect -483 -250 -477 -246
rect -402 -247 -396 -243
rect -402 -249 -392 -247
rect -487 -251 -477 -250
rect -402 -252 -392 -251
rect -587 -261 -571 -257
rect -487 -254 -477 -253
rect -487 -258 -481 -254
rect -398 -256 -392 -252
rect -591 -262 -571 -261
rect -591 -271 -571 -264
rect -591 -274 -571 -273
rect -591 -278 -575 -274
rect -487 -276 -471 -272
rect -491 -277 -471 -276
rect -491 -280 -471 -279
rect -491 -284 -475 -280
rect -583 -288 -577 -284
rect -587 -289 -577 -288
rect -587 -292 -577 -291
rect -587 -296 -581 -292
rect -487 -300 -471 -296
rect -491 -301 -471 -300
rect -491 -304 -471 -303
rect -491 -308 -475 -304
rect -587 -314 -571 -310
rect -591 -315 -571 -314
rect -591 -318 -571 -317
rect -591 -322 -575 -318
rect -304 -282 -299 -266
rect -300 -286 -299 -282
rect -297 -286 -289 -266
rect -287 -270 -286 -266
rect 61 -199 77 -195
rect 57 -200 77 -199
rect 57 -203 77 -202
rect 57 -207 73 -203
rect -287 -286 -282 -270
rect 61 -223 77 -219
rect 57 -224 77 -223
rect 57 -227 77 -226
rect 57 -231 73 -227
rect -105 -259 -100 -253
rect -101 -263 -100 -259
rect -98 -257 -96 -253
rect -92 -257 -90 -253
rect -98 -263 -90 -257
rect -88 -259 -83 -253
rect -54 -255 -49 -239
rect -50 -259 -49 -255
rect -47 -259 -39 -239
rect -37 -243 -36 -239
rect -37 -259 -32 -243
rect -23 -245 -18 -239
rect -19 -249 -18 -245
rect -16 -243 -15 -239
rect -16 -249 -11 -243
rect -88 -263 -87 -259
rect -261 -292 -256 -286
rect -257 -296 -256 -292
rect -254 -290 -252 -286
rect -248 -290 -246 -286
rect -254 -296 -246 -290
rect -244 -292 -239 -286
rect -233 -288 -228 -282
rect -229 -292 -228 -288
rect -226 -286 -225 -282
rect -226 -292 -221 -286
rect -244 -296 -243 -292
rect -414 -324 -413 -320
rect -418 -330 -413 -324
rect -411 -326 -406 -320
rect -411 -330 -410 -326
rect -393 -324 -392 -320
rect -587 -338 -571 -334
rect -591 -339 -571 -338
rect -397 -340 -392 -324
rect -390 -340 -382 -320
rect -380 -336 -375 -320
rect 6 -319 7 -315
rect -380 -340 -379 -336
rect -346 -340 -341 -334
rect -591 -342 -571 -341
rect -591 -346 -575 -342
rect -342 -344 -341 -340
rect -339 -338 -337 -334
rect -333 -338 -331 -334
rect -339 -344 -331 -338
rect -329 -340 -324 -334
rect -329 -344 -328 -340
rect 2 -325 7 -319
rect 9 -321 14 -315
rect 9 -325 10 -321
rect 20 -325 25 -319
rect 24 -329 25 -325
rect 27 -323 29 -319
rect 33 -323 35 -319
rect 27 -329 35 -323
rect 37 -325 42 -319
rect 37 -329 38 -325
rect -539 -385 -534 -379
rect -535 -389 -534 -385
rect -532 -383 -531 -379
rect -532 -389 -527 -383
rect -275 -361 -274 -357
rect -279 -367 -274 -361
rect -272 -361 -270 -357
rect -266 -361 -265 -357
rect -272 -367 -265 -361
rect -263 -363 -258 -357
rect -263 -367 -262 -363
rect -242 -362 -237 -356
rect -238 -366 -237 -362
rect -235 -362 -230 -356
rect -235 -366 -234 -362
rect 54 -335 59 -319
rect 58 -339 59 -335
rect 61 -339 69 -319
rect 71 -323 72 -319
rect 71 -339 76 -323
rect 85 -325 90 -319
rect 89 -329 90 -325
rect 92 -323 93 -319
rect 92 -329 97 -323
rect 120 -335 125 -329
rect 124 -339 125 -335
rect 127 -333 129 -329
rect 133 -333 135 -329
rect 127 -339 135 -333
rect 137 -335 142 -329
rect 148 -331 153 -325
rect 152 -335 153 -331
rect 155 -329 156 -325
rect 155 -335 160 -329
rect 137 -339 138 -335
rect 179 -347 184 -331
rect 183 -351 184 -347
rect 186 -351 194 -331
rect 196 -335 197 -331
rect 196 -351 201 -335
rect -515 -411 -510 -405
rect -511 -415 -510 -411
rect -508 -409 -506 -405
rect -502 -409 -500 -405
rect -508 -415 -500 -409
rect -498 -411 -493 -405
rect -487 -407 -482 -401
rect -483 -411 -482 -407
rect -480 -405 -479 -401
rect -480 -411 -475 -405
rect -193 -377 -192 -373
rect -197 -383 -192 -377
rect -190 -379 -185 -373
rect -190 -383 -189 -379
rect -172 -377 -171 -373
rect -176 -393 -171 -377
rect -169 -393 -161 -373
rect -159 -389 -154 -373
rect 159 -367 165 -363
rect 159 -368 169 -367
rect 159 -372 169 -370
rect 163 -376 169 -372
rect 159 -378 169 -376
rect 159 -381 169 -380
rect 159 -385 165 -381
rect -159 -393 -158 -389
rect -498 -415 -497 -411
rect -606 -425 -605 -421
rect -610 -431 -605 -425
rect -603 -425 -601 -421
rect -597 -425 -596 -421
rect -603 -431 -596 -425
rect -594 -427 -589 -421
rect -594 -431 -593 -427
rect -573 -426 -568 -420
rect -569 -430 -568 -426
rect -566 -426 -561 -420
rect -566 -430 -565 -426
rect -466 -423 -461 -407
rect -462 -427 -461 -423
rect -459 -427 -451 -407
rect -449 -411 -448 -407
rect -139 -394 -134 -388
rect -135 -398 -134 -394
rect -132 -392 -130 -388
rect -126 -392 -124 -388
rect -132 -398 -124 -392
rect -122 -394 -117 -388
rect -122 -398 -121 -394
rect -84 -404 -79 -398
rect -80 -408 -79 -404
rect -77 -404 -72 -398
rect -77 -408 -76 -404
rect -56 -405 -51 -399
rect -449 -427 -444 -411
rect -412 -413 -411 -409
rect -416 -419 -411 -413
rect -409 -413 -407 -409
rect -403 -413 -402 -409
rect -409 -419 -402 -413
rect -400 -415 -395 -409
rect -400 -419 -399 -415
rect -379 -414 -374 -408
rect -375 -418 -374 -414
rect -372 -414 -367 -408
rect -52 -409 -51 -405
rect -49 -403 -48 -399
rect -44 -403 -42 -399
rect -49 -409 -42 -403
rect -40 -403 -39 -399
rect -40 -409 -35 -403
rect -372 -418 -371 -414
rect -564 -458 -559 -452
rect -560 -462 -559 -458
rect -557 -458 -550 -452
rect -557 -462 -555 -458
rect -551 -462 -550 -458
rect -548 -456 -547 -452
rect -496 -452 -495 -448
rect -548 -462 -543 -456
rect -523 -457 -522 -453
rect -527 -463 -522 -457
rect -520 -457 -519 -453
rect -520 -463 -515 -457
rect -500 -458 -495 -452
rect -493 -454 -485 -448
rect -493 -458 -491 -454
rect -487 -458 -485 -454
rect -483 -452 -482 -448
rect -483 -458 -478 -452
rect -462 -453 -461 -449
rect -466 -469 -461 -453
rect -459 -469 -451 -449
rect -449 -465 -444 -449
rect -404 -458 -399 -452
rect -400 -462 -399 -458
rect -397 -458 -390 -452
rect -397 -462 -395 -458
rect -391 -462 -390 -458
rect -388 -456 -387 -452
rect -336 -452 -335 -448
rect -388 -462 -383 -456
rect -363 -457 -362 -453
rect -449 -469 -448 -465
rect -367 -463 -362 -457
rect -360 -457 -359 -453
rect -360 -463 -355 -457
rect -340 -458 -335 -452
rect -333 -454 -325 -448
rect -333 -458 -331 -454
rect -327 -458 -325 -454
rect -323 -452 -322 -448
rect -323 -458 -318 -452
rect -302 -453 -301 -449
rect -306 -469 -301 -453
rect -299 -469 -291 -449
rect -289 -465 -284 -449
rect -255 -455 -250 -449
rect -251 -459 -250 -455
rect -248 -455 -241 -449
rect -248 -459 -246 -455
rect -242 -459 -241 -455
rect -239 -453 -238 -449
rect -187 -449 -186 -445
rect -239 -459 -234 -453
rect -214 -454 -213 -450
rect -289 -469 -288 -465
rect -218 -460 -213 -454
rect -211 -454 -210 -450
rect -211 -460 -206 -454
rect -191 -455 -186 -449
rect -184 -451 -176 -445
rect -184 -455 -182 -451
rect -178 -455 -176 -451
rect -174 -449 -173 -445
rect -174 -455 -169 -449
rect -153 -450 -152 -446
rect -157 -466 -152 -450
rect -150 -466 -142 -446
rect -140 -462 -135 -446
rect -103 -455 -98 -449
rect -99 -459 -98 -455
rect -96 -455 -89 -449
rect -96 -459 -94 -455
rect -90 -459 -89 -455
rect -87 -453 -86 -449
rect -35 -449 -34 -445
rect -87 -459 -82 -453
rect -62 -454 -61 -450
rect -140 -466 -139 -462
rect -66 -460 -61 -454
rect -59 -454 -58 -450
rect -59 -460 -54 -454
rect -39 -455 -34 -449
rect -32 -451 -24 -445
rect -32 -455 -30 -451
rect -26 -455 -24 -451
rect -22 -449 -21 -445
rect -22 -455 -17 -449
rect -1 -450 0 -446
rect -5 -466 0 -450
rect 2 -466 10 -446
rect 12 -462 17 -446
rect 12 -466 13 -462
rect 49 -460 54 -444
rect 53 -464 54 -460
rect 56 -464 64 -444
rect 66 -448 67 -444
rect 66 -464 71 -448
rect 83 -460 88 -444
rect 87 -464 88 -460
rect 90 -464 98 -444
rect 100 -448 101 -444
rect 100 -464 105 -448
rect -568 -548 -562 -544
rect -572 -549 -562 -548
rect -489 -549 -483 -545
rect -407 -546 -401 -542
rect -411 -547 -401 -546
rect -323 -547 -317 -543
rect -241 -546 -235 -542
rect -245 -547 -235 -546
rect -155 -546 -149 -542
rect -159 -547 -149 -546
rect -327 -548 -317 -547
rect -493 -550 -483 -549
rect -572 -552 -562 -551
rect -572 -556 -566 -552
rect -493 -553 -483 -552
rect -493 -557 -487 -553
rect -411 -550 -401 -549
rect -70 -547 -64 -543
rect -74 -548 -64 -547
rect 13 -547 19 -543
rect 9 -548 19 -547
rect 97 -547 103 -543
rect 93 -548 103 -547
rect -411 -554 -405 -550
rect -327 -551 -317 -550
rect -327 -555 -321 -551
rect -245 -550 -235 -549
rect -245 -554 -239 -550
rect -159 -550 -149 -549
rect -159 -554 -153 -550
rect -74 -551 -64 -550
rect -74 -555 -68 -551
rect 9 -551 19 -550
rect 9 -555 15 -551
rect 93 -551 103 -550
rect 93 -555 99 -551
rect -572 -564 -556 -560
rect -576 -565 -556 -564
rect -493 -565 -477 -561
rect -411 -562 -395 -558
rect -415 -563 -395 -562
rect -327 -563 -311 -559
rect -245 -562 -229 -558
rect -249 -563 -229 -562
rect -159 -562 -143 -558
rect -163 -563 -143 -562
rect -74 -563 -58 -559
rect -331 -564 -311 -563
rect -497 -566 -477 -565
rect -576 -574 -556 -567
rect -497 -575 -477 -568
rect -415 -572 -395 -565
rect -78 -564 -58 -563
rect 9 -563 25 -559
rect 5 -564 25 -563
rect 93 -563 109 -559
rect 89 -564 109 -563
rect -331 -573 -311 -566
rect -249 -572 -229 -565
rect -163 -572 -143 -565
rect -576 -577 -556 -576
rect -576 -581 -560 -577
rect -497 -578 -477 -577
rect -497 -582 -481 -578
rect -415 -575 -395 -574
rect -78 -573 -58 -566
rect 5 -573 25 -566
rect 89 -573 109 -566
rect -415 -579 -399 -575
rect -331 -576 -311 -575
rect -331 -580 -315 -576
rect -249 -575 -229 -574
rect -249 -579 -233 -575
rect -163 -575 -143 -574
rect -163 -579 -147 -575
rect -78 -576 -58 -575
rect -78 -580 -62 -576
rect 5 -576 25 -575
rect 5 -580 21 -576
rect 89 -576 109 -575
rect 89 -580 105 -576
rect -572 -589 -556 -585
rect -576 -590 -556 -589
rect -493 -590 -477 -586
rect -411 -587 -395 -583
rect -415 -588 -395 -587
rect -327 -588 -311 -584
rect -245 -587 -229 -583
rect -249 -588 -229 -587
rect -159 -587 -143 -583
rect -163 -588 -143 -587
rect -74 -588 -58 -584
rect -331 -589 -311 -588
rect -497 -591 -477 -590
rect -576 -599 -556 -592
rect -497 -600 -477 -593
rect -415 -597 -395 -590
rect -78 -589 -58 -588
rect 9 -588 25 -584
rect 5 -589 25 -588
rect 93 -588 109 -584
rect 89 -589 109 -588
rect -331 -598 -311 -591
rect -249 -597 -229 -590
rect -163 -597 -143 -590
rect -576 -602 -556 -601
rect -576 -606 -560 -602
rect -497 -603 -477 -602
rect -497 -607 -481 -603
rect -415 -600 -395 -599
rect -78 -598 -58 -591
rect 5 -598 25 -591
rect 89 -598 109 -591
rect -415 -604 -399 -600
rect -331 -601 -311 -600
rect -331 -605 -315 -601
rect -249 -600 -229 -599
rect -249 -604 -233 -600
rect -163 -600 -143 -599
rect -163 -604 -147 -600
rect -78 -601 -58 -600
rect -78 -605 -62 -601
rect 5 -601 25 -600
rect 5 -605 21 -601
rect 89 -601 109 -600
rect 89 -605 105 -601
rect -568 -616 -562 -612
rect -572 -617 -562 -616
rect -489 -617 -483 -613
rect -407 -614 -401 -610
rect -411 -615 -401 -614
rect -323 -615 -317 -611
rect -241 -614 -235 -610
rect -245 -615 -235 -614
rect -155 -614 -149 -610
rect -159 -615 -149 -614
rect -327 -616 -317 -615
rect -493 -618 -483 -617
rect -572 -620 -562 -619
rect -572 -624 -566 -620
rect -493 -621 -483 -620
rect -493 -625 -487 -621
rect -411 -618 -401 -617
rect -70 -615 -64 -611
rect -74 -616 -64 -615
rect 13 -615 19 -611
rect 9 -616 19 -615
rect 97 -615 103 -611
rect 93 -616 103 -615
rect -411 -622 -405 -618
rect -327 -619 -317 -618
rect -327 -623 -321 -619
rect -245 -618 -235 -617
rect -245 -622 -239 -618
rect -159 -618 -149 -617
rect -159 -622 -153 -618
rect -74 -619 -64 -618
rect -74 -623 -68 -619
rect 9 -619 19 -618
rect 9 -623 15 -619
rect 93 -619 103 -618
rect 93 -623 99 -619
rect -572 -642 -556 -638
rect -576 -643 -556 -642
rect -493 -643 -477 -639
rect -411 -640 -395 -636
rect -415 -641 -395 -640
rect -327 -641 -311 -637
rect -245 -640 -229 -636
rect -249 -641 -229 -640
rect -159 -640 -143 -636
rect -163 -641 -143 -640
rect -331 -642 -311 -641
rect -497 -644 -477 -643
rect -576 -646 -556 -645
rect -576 -650 -560 -646
rect -497 -647 -477 -646
rect -497 -651 -481 -647
rect -415 -644 -395 -643
rect -74 -641 -58 -637
rect -78 -642 -58 -641
rect 9 -641 25 -637
rect 5 -642 25 -641
rect 93 -641 109 -637
rect 89 -642 109 -641
rect -415 -648 -399 -644
rect -331 -645 -311 -644
rect -331 -649 -315 -645
rect -249 -644 -229 -643
rect -249 -648 -233 -644
rect -163 -644 -143 -643
rect -163 -648 -147 -644
rect -78 -645 -58 -644
rect -78 -649 -62 -645
rect 5 -645 25 -644
rect 5 -649 21 -645
rect 89 -645 109 -644
rect 89 -649 105 -645
rect -572 -666 -556 -662
rect -576 -667 -556 -666
rect -493 -667 -477 -663
rect -411 -664 -395 -660
rect -415 -665 -395 -664
rect -327 -665 -311 -661
rect -245 -664 -229 -660
rect -249 -665 -229 -664
rect -159 -664 -143 -660
rect -163 -665 -143 -664
rect -331 -666 -311 -665
rect -497 -668 -477 -667
rect -576 -670 -556 -669
rect -576 -674 -560 -670
rect -497 -671 -477 -670
rect -497 -675 -481 -671
rect -415 -668 -395 -667
rect -74 -665 -58 -661
rect -78 -666 -58 -665
rect 9 -665 25 -661
rect 5 -666 25 -665
rect 93 -665 109 -661
rect 89 -666 109 -665
rect -415 -672 -399 -668
rect -331 -669 -311 -668
rect -331 -673 -315 -669
rect -249 -668 -229 -667
rect -249 -672 -233 -668
rect -163 -668 -143 -667
rect -163 -672 -147 -668
rect -78 -669 -58 -668
rect -78 -673 -62 -669
rect 5 -669 25 -668
rect 5 -673 21 -669
rect 89 -669 109 -668
rect 89 -673 105 -669
<< pdiffusion >>
rect -118 50 -102 54
rect -118 49 -98 50
rect -118 46 -98 47
rect -114 42 -98 46
rect -118 26 -102 30
rect -118 25 -98 26
rect -118 22 -98 23
rect -114 18 -98 22
rect -118 1 -102 5
rect -118 0 -98 1
rect -118 -3 -98 -2
rect -114 -7 -98 -3
rect -118 -24 -102 -20
rect -118 -25 -98 -24
rect -118 -28 -98 -27
rect -114 -32 -98 -28
rect -321 -38 -305 -34
rect -321 -39 -301 -38
rect -321 -42 -301 -41
rect -317 -46 -301 -42
rect -118 -42 -102 -38
rect -118 -43 -98 -42
rect -118 -46 -98 -45
rect -114 -50 -98 -46
rect -321 -62 -305 -58
rect -321 -63 -301 -62
rect -118 -60 -102 -56
rect -118 -61 -98 -60
rect -321 -66 -301 -65
rect -317 -70 -301 -66
rect -118 -69 -98 -63
rect -118 -72 -98 -71
rect -114 -76 -98 -72
rect -321 -87 -305 -83
rect -321 -88 -301 -87
rect -118 -84 -102 -80
rect 25 -81 41 -77
rect 25 -82 45 -81
rect -118 -85 -98 -84
rect 25 -85 45 -84
rect -321 -91 -301 -90
rect -317 -95 -301 -91
rect -118 -93 -98 -87
rect 29 -89 45 -85
rect -118 -96 -98 -95
rect -114 -100 -98 -96
rect 25 -105 41 -101
rect 25 -106 45 -105
rect -321 -112 -305 -108
rect -321 -113 -301 -112
rect 25 -109 45 -108
rect 29 -113 45 -109
rect -321 -116 -301 -115
rect -317 -120 -301 -116
rect -321 -130 -305 -126
rect -321 -131 -301 -130
rect 25 -130 41 -126
rect 25 -131 45 -130
rect -321 -134 -301 -133
rect -317 -138 -301 -134
rect 25 -134 45 -133
rect -73 -139 -57 -135
rect -73 -140 -53 -139
rect 29 -138 45 -134
rect -73 -143 -53 -142
rect -321 -148 -305 -144
rect -69 -147 -53 -143
rect -321 -149 -301 -148
rect -523 -158 -507 -154
rect -523 -159 -503 -158
rect -321 -157 -301 -151
rect -321 -160 -301 -159
rect -523 -162 -503 -161
rect -519 -166 -503 -162
rect -317 -164 -301 -160
rect -321 -172 -305 -168
rect -321 -173 -301 -172
rect -523 -182 -507 -178
rect -523 -183 -503 -182
rect -321 -181 -301 -175
rect -321 -184 -301 -183
rect -523 -186 -503 -185
rect -519 -190 -503 -186
rect -317 -188 -301 -184
rect -208 -185 -203 -169
rect -204 -189 -203 -185
rect -201 -173 -200 -169
rect -201 -189 -196 -173
rect -190 -183 -185 -147
rect -186 -187 -185 -183
rect -183 -187 -175 -147
rect -173 -151 -172 -147
rect -173 -187 -168 -151
rect -143 -151 -142 -147
rect -147 -167 -142 -151
rect -140 -163 -132 -147
rect -140 -167 -138 -163
rect -134 -167 -132 -163
rect -130 -151 -129 -147
rect -130 -167 -125 -151
rect -95 -157 -59 -153
rect -95 -158 -55 -157
rect 25 -155 41 -151
rect 25 -156 45 -155
rect 25 -159 45 -158
rect -95 -168 -55 -160
rect 29 -163 45 -159
rect -95 -171 -55 -170
rect -91 -175 -55 -171
rect 25 -173 41 -169
rect 25 -174 45 -173
rect 25 -177 45 -176
rect 29 -181 45 -177
rect -623 -196 -607 -192
rect -623 -197 -603 -196
rect -623 -200 -603 -199
rect -619 -204 -603 -200
rect -523 -207 -507 -203
rect -523 -208 -503 -207
rect -523 -211 -503 -210
rect -519 -215 -503 -211
rect 25 -191 41 -187
rect 25 -192 45 -191
rect -101 -199 -100 -195
rect -623 -220 -607 -216
rect -623 -221 -603 -220
rect -372 -220 -356 -216
rect -376 -221 -356 -220
rect -623 -224 -603 -223
rect -619 -228 -603 -224
rect -523 -232 -507 -228
rect -523 -233 -503 -232
rect -376 -224 -356 -223
rect -376 -228 -360 -224
rect -300 -232 -299 -228
rect -523 -236 -503 -235
rect -623 -245 -607 -241
rect -623 -246 -603 -245
rect -519 -240 -503 -236
rect -370 -238 -334 -234
rect -374 -239 -334 -238
rect -623 -249 -603 -248
rect -619 -253 -603 -249
rect -523 -250 -507 -246
rect -523 -251 -503 -250
rect -374 -249 -334 -241
rect -304 -248 -299 -232
rect -297 -244 -289 -228
rect -297 -248 -295 -244
rect -291 -248 -289 -244
rect -287 -232 -286 -228
rect -287 -248 -282 -232
rect -257 -232 -256 -228
rect -523 -254 -503 -253
rect -519 -258 -503 -254
rect -374 -252 -334 -251
rect -374 -256 -338 -252
rect -623 -270 -607 -266
rect -623 -271 -603 -270
rect -523 -268 -507 -264
rect -523 -269 -503 -268
rect -623 -274 -603 -273
rect -619 -278 -603 -274
rect -523 -277 -503 -271
rect -523 -280 -503 -279
rect -519 -284 -503 -280
rect -623 -288 -607 -284
rect -623 -289 -603 -288
rect -393 -286 -392 -282
rect -623 -292 -603 -291
rect -619 -296 -603 -292
rect -523 -292 -507 -288
rect -523 -293 -503 -292
rect -523 -301 -503 -295
rect -623 -306 -607 -302
rect -623 -307 -603 -306
rect -523 -304 -503 -303
rect -519 -308 -503 -304
rect -418 -304 -413 -288
rect -414 -308 -413 -304
rect -411 -292 -410 -288
rect -411 -308 -406 -292
rect -397 -302 -392 -286
rect -390 -298 -382 -282
rect -390 -302 -388 -298
rect -384 -302 -382 -298
rect -380 -286 -379 -282
rect -380 -302 -375 -286
rect -623 -315 -603 -309
rect -623 -318 -603 -317
rect -619 -322 -603 -318
rect -346 -312 -341 -276
rect -342 -316 -341 -312
rect -339 -316 -331 -276
rect -329 -280 -328 -276
rect -329 -316 -324 -280
rect -261 -268 -256 -232
rect -254 -268 -246 -228
rect -244 -264 -239 -228
rect -105 -235 -100 -199
rect -98 -235 -90 -195
rect -88 -231 -83 -195
rect 25 -200 45 -194
rect -50 -205 -49 -201
rect -54 -221 -49 -205
rect -47 -217 -39 -201
rect -47 -221 -45 -217
rect -41 -221 -39 -217
rect -37 -205 -36 -201
rect 25 -203 45 -202
rect -37 -221 -32 -205
rect 29 -207 45 -203
rect -19 -211 -18 -207
rect -88 -235 -87 -231
rect -244 -268 -243 -264
rect -229 -254 -228 -250
rect -233 -270 -228 -254
rect -226 -266 -221 -250
rect -23 -227 -18 -211
rect -16 -223 -11 -207
rect 25 -215 41 -211
rect 25 -216 45 -215
rect -16 -227 -15 -223
rect 25 -224 45 -218
rect 25 -227 45 -226
rect 29 -231 45 -227
rect -226 -270 -225 -266
rect 2 -299 7 -283
rect 6 -303 7 -299
rect 9 -287 10 -283
rect 9 -303 14 -287
rect 20 -297 25 -261
rect 24 -301 25 -297
rect 27 -301 35 -261
rect 37 -265 38 -261
rect 37 -301 42 -265
rect 124 -275 125 -271
rect 58 -285 59 -281
rect 54 -301 59 -285
rect 61 -297 69 -281
rect 61 -301 63 -297
rect 67 -301 69 -297
rect 71 -285 72 -281
rect 71 -301 76 -285
rect 89 -291 90 -287
rect -623 -330 -607 -326
rect -623 -331 -603 -330
rect -623 -339 -603 -333
rect -623 -342 -603 -341
rect -619 -346 -603 -342
rect -279 -340 -274 -324
rect -275 -344 -274 -340
rect -272 -338 -265 -324
rect -272 -342 -270 -338
rect -266 -342 -265 -338
rect -272 -344 -265 -342
rect -263 -328 -262 -324
rect -263 -344 -258 -328
rect -238 -328 -237 -324
rect -242 -344 -237 -328
rect -235 -340 -230 -324
rect 85 -307 90 -291
rect 92 -303 97 -287
rect 92 -307 93 -303
rect 120 -311 125 -275
rect 127 -311 135 -271
rect 137 -307 142 -271
rect 137 -311 138 -307
rect 152 -297 153 -293
rect -235 -344 -234 -340
rect -172 -339 -171 -335
rect -535 -351 -534 -347
rect -539 -367 -534 -351
rect -532 -363 -527 -347
rect -532 -367 -531 -363
rect -511 -351 -510 -347
rect -610 -404 -605 -388
rect -606 -408 -605 -404
rect -603 -402 -596 -388
rect -603 -406 -601 -402
rect -597 -406 -596 -402
rect -603 -408 -596 -406
rect -594 -392 -593 -388
rect -594 -408 -589 -392
rect -569 -392 -568 -388
rect -573 -408 -568 -392
rect -566 -404 -561 -388
rect -515 -387 -510 -351
rect -508 -387 -500 -347
rect -498 -383 -493 -347
rect -498 -387 -497 -383
rect -483 -373 -482 -369
rect -566 -408 -565 -404
rect -487 -389 -482 -373
rect -480 -385 -475 -369
rect -480 -389 -479 -385
rect -462 -373 -461 -369
rect -466 -389 -461 -373
rect -459 -385 -451 -369
rect -459 -389 -457 -385
rect -453 -389 -451 -385
rect -449 -373 -448 -369
rect -449 -389 -444 -373
rect -197 -357 -192 -341
rect -193 -361 -192 -357
rect -190 -345 -189 -341
rect -190 -361 -185 -345
rect -176 -355 -171 -339
rect -169 -351 -161 -335
rect -169 -355 -167 -351
rect -163 -355 -161 -351
rect -159 -339 -158 -335
rect -159 -355 -154 -339
rect -139 -366 -134 -330
rect -135 -370 -134 -366
rect -132 -370 -124 -330
rect -122 -334 -121 -330
rect -122 -370 -117 -334
rect 148 -313 153 -297
rect 155 -309 160 -293
rect 155 -313 156 -309
rect 183 -297 184 -293
rect 179 -313 184 -297
rect 186 -309 194 -293
rect 186 -313 188 -309
rect 192 -313 194 -309
rect 196 -297 197 -293
rect 196 -313 201 -297
rect -416 -392 -411 -376
rect -412 -396 -411 -392
rect -409 -390 -402 -376
rect -409 -394 -407 -390
rect -403 -394 -402 -390
rect -409 -396 -402 -394
rect -400 -380 -399 -376
rect -400 -396 -395 -380
rect -375 -380 -374 -376
rect -379 -396 -374 -380
rect -372 -392 -367 -376
rect -372 -396 -371 -392
rect -84 -382 -79 -366
rect -80 -386 -79 -382
rect -77 -370 -76 -366
rect -77 -386 -72 -370
rect -52 -370 -51 -366
rect -56 -386 -51 -370
rect -49 -380 -42 -366
rect -49 -384 -48 -380
rect -44 -384 -42 -380
rect -49 -386 -42 -384
rect -40 -382 -35 -366
rect 105 -367 141 -363
rect 101 -368 141 -367
rect 101 -378 141 -370
rect -40 -386 -39 -382
rect 101 -381 141 -380
rect 101 -385 137 -381
rect 53 -410 54 -406
rect 49 -426 54 -410
rect 56 -422 64 -406
rect 56 -426 58 -422
rect 62 -426 64 -422
rect 66 -410 67 -406
rect 66 -426 71 -410
rect 87 -410 88 -406
rect 83 -426 88 -410
rect 90 -422 98 -406
rect 90 -426 92 -422
rect 96 -426 98 -422
rect 100 -410 101 -406
rect 100 -426 105 -410
rect -560 -479 -559 -475
rect -564 -495 -559 -479
rect -557 -477 -550 -475
rect -557 -481 -555 -477
rect -551 -481 -550 -477
rect -557 -495 -550 -481
rect -548 -491 -543 -475
rect -548 -495 -547 -491
rect -527 -491 -522 -475
rect -523 -495 -522 -491
rect -520 -479 -519 -475
rect -520 -495 -515 -479
rect -500 -512 -495 -476
rect -496 -516 -495 -512
rect -493 -516 -485 -476
rect -483 -480 -482 -476
rect -483 -516 -478 -480
rect -400 -479 -399 -475
rect -466 -503 -461 -487
rect -462 -507 -461 -503
rect -459 -491 -457 -487
rect -453 -491 -451 -487
rect -459 -507 -451 -491
rect -449 -503 -444 -487
rect -404 -495 -399 -479
rect -397 -477 -390 -475
rect -397 -481 -395 -477
rect -391 -481 -390 -477
rect -397 -495 -390 -481
rect -388 -491 -383 -475
rect -388 -495 -387 -491
rect -367 -491 -362 -475
rect -363 -495 -362 -491
rect -360 -479 -359 -475
rect -360 -495 -355 -479
rect -449 -507 -448 -503
rect -340 -512 -335 -476
rect -336 -516 -335 -512
rect -333 -516 -325 -476
rect -323 -480 -322 -476
rect -323 -516 -318 -480
rect -251 -476 -250 -472
rect -306 -503 -301 -487
rect -302 -507 -301 -503
rect -299 -491 -297 -487
rect -293 -491 -291 -487
rect -299 -507 -291 -491
rect -289 -503 -284 -487
rect -255 -492 -250 -476
rect -248 -474 -241 -472
rect -248 -478 -246 -474
rect -242 -478 -241 -474
rect -248 -492 -241 -478
rect -239 -488 -234 -472
rect -239 -492 -238 -488
rect -218 -488 -213 -472
rect -214 -492 -213 -488
rect -211 -476 -210 -472
rect -211 -492 -206 -476
rect -289 -507 -288 -503
rect -191 -509 -186 -473
rect -187 -513 -186 -509
rect -184 -513 -176 -473
rect -174 -477 -173 -473
rect -174 -513 -169 -477
rect -99 -476 -98 -472
rect -157 -500 -152 -484
rect -153 -504 -152 -500
rect -150 -488 -148 -484
rect -144 -488 -142 -484
rect -150 -504 -142 -488
rect -140 -500 -135 -484
rect -103 -492 -98 -476
rect -96 -474 -89 -472
rect -96 -478 -94 -474
rect -90 -478 -89 -474
rect -96 -492 -89 -478
rect -87 -488 -82 -472
rect -87 -492 -86 -488
rect -66 -488 -61 -472
rect -62 -492 -61 -488
rect -59 -476 -58 -472
rect -59 -492 -54 -476
rect -140 -504 -139 -500
rect -39 -509 -34 -473
rect -35 -513 -34 -509
rect -32 -513 -24 -473
rect -22 -477 -21 -473
rect -22 -513 -17 -477
rect -5 -500 0 -484
rect -1 -504 0 -500
rect 2 -488 4 -484
rect 8 -488 10 -484
rect 2 -504 10 -488
rect 12 -500 17 -484
rect 12 -504 13 -500
rect -608 -548 -592 -544
rect -608 -549 -588 -548
rect -529 -549 -513 -545
rect -529 -550 -509 -549
rect -447 -546 -431 -542
rect -447 -547 -427 -546
rect -363 -547 -347 -543
rect -363 -548 -343 -547
rect -281 -546 -265 -542
rect -281 -547 -261 -546
rect -195 -546 -179 -542
rect -195 -547 -175 -546
rect -110 -547 -94 -543
rect -447 -550 -427 -549
rect -608 -552 -588 -551
rect -604 -556 -588 -552
rect -529 -553 -509 -552
rect -525 -557 -509 -553
rect -443 -554 -427 -550
rect -110 -548 -90 -547
rect -27 -547 -11 -543
rect -27 -548 -7 -547
rect 57 -547 73 -543
rect 57 -548 77 -547
rect -281 -550 -261 -549
rect -363 -551 -343 -550
rect -359 -555 -343 -551
rect -277 -554 -261 -550
rect -195 -550 -175 -549
rect -191 -554 -175 -550
rect -110 -551 -90 -550
rect -106 -555 -90 -551
rect -27 -551 -7 -550
rect -23 -555 -7 -551
rect 57 -551 77 -550
rect 61 -555 77 -551
rect -608 -573 -592 -569
rect -608 -574 -588 -573
rect -529 -574 -513 -570
rect -529 -575 -509 -574
rect -447 -571 -431 -567
rect -447 -572 -427 -571
rect -363 -572 -347 -568
rect -363 -573 -343 -572
rect -281 -571 -265 -567
rect -281 -572 -261 -571
rect -195 -571 -179 -567
rect -195 -572 -175 -571
rect -110 -572 -94 -568
rect -447 -575 -427 -574
rect -608 -577 -588 -576
rect -604 -581 -588 -577
rect -529 -578 -509 -577
rect -525 -582 -509 -578
rect -443 -579 -427 -575
rect -110 -573 -90 -572
rect -27 -572 -11 -568
rect -27 -573 -7 -572
rect 57 -572 73 -568
rect 57 -573 77 -572
rect -281 -575 -261 -574
rect -363 -576 -343 -575
rect -359 -580 -343 -576
rect -277 -579 -261 -575
rect -195 -575 -175 -574
rect -191 -579 -175 -575
rect -110 -576 -90 -575
rect -106 -580 -90 -576
rect -27 -576 -7 -575
rect -23 -580 -7 -576
rect 57 -576 77 -575
rect 61 -580 77 -576
rect -608 -598 -592 -594
rect -608 -599 -588 -598
rect -529 -599 -513 -595
rect -529 -600 -509 -599
rect -447 -596 -431 -592
rect -447 -597 -427 -596
rect -363 -597 -347 -593
rect -363 -598 -343 -597
rect -281 -596 -265 -592
rect -281 -597 -261 -596
rect -195 -596 -179 -592
rect -195 -597 -175 -596
rect -110 -597 -94 -593
rect -447 -600 -427 -599
rect -608 -602 -588 -601
rect -604 -606 -588 -602
rect -529 -603 -509 -602
rect -525 -607 -509 -603
rect -443 -604 -427 -600
rect -110 -598 -90 -597
rect -27 -597 -11 -593
rect -27 -598 -7 -597
rect 57 -597 73 -593
rect 57 -598 77 -597
rect -281 -600 -261 -599
rect -363 -601 -343 -600
rect -359 -605 -343 -601
rect -277 -604 -261 -600
rect -195 -600 -175 -599
rect -191 -604 -175 -600
rect -110 -601 -90 -600
rect -106 -605 -90 -601
rect -27 -601 -7 -600
rect -23 -605 -7 -601
rect 57 -601 77 -600
rect 61 -605 77 -601
rect -608 -616 -592 -612
rect -608 -617 -588 -616
rect -529 -617 -513 -613
rect -529 -618 -509 -617
rect -447 -614 -431 -610
rect -447 -615 -427 -614
rect -363 -615 -347 -611
rect -363 -616 -343 -615
rect -281 -614 -265 -610
rect -281 -615 -261 -614
rect -195 -614 -179 -610
rect -195 -615 -175 -614
rect -110 -615 -94 -611
rect -447 -618 -427 -617
rect -608 -620 -588 -619
rect -604 -624 -588 -620
rect -529 -621 -509 -620
rect -525 -625 -509 -621
rect -443 -622 -427 -618
rect -110 -616 -90 -615
rect -27 -615 -11 -611
rect -27 -616 -7 -615
rect 57 -615 73 -611
rect 57 -616 77 -615
rect -281 -618 -261 -617
rect -363 -619 -343 -618
rect -359 -623 -343 -619
rect -277 -622 -261 -618
rect -195 -618 -175 -617
rect -191 -622 -175 -618
rect -110 -619 -90 -618
rect -106 -623 -90 -619
rect -27 -619 -7 -618
rect -23 -623 -7 -619
rect 57 -619 77 -618
rect 61 -623 77 -619
rect -608 -634 -592 -630
rect -608 -635 -588 -634
rect -529 -635 -513 -631
rect -447 -632 -431 -628
rect -447 -633 -427 -632
rect -363 -633 -347 -629
rect -281 -632 -265 -628
rect -281 -633 -261 -632
rect -195 -632 -179 -628
rect -195 -633 -175 -632
rect -110 -633 -94 -629
rect -363 -634 -343 -633
rect -529 -636 -509 -635
rect -608 -643 -588 -637
rect -529 -644 -509 -638
rect -447 -641 -427 -635
rect -110 -634 -90 -633
rect -27 -633 -11 -629
rect -27 -634 -7 -633
rect 57 -633 73 -629
rect 57 -634 77 -633
rect -363 -642 -343 -636
rect -281 -641 -261 -635
rect -195 -641 -175 -635
rect -447 -644 -427 -643
rect -608 -646 -588 -645
rect -604 -650 -588 -646
rect -529 -647 -509 -646
rect -525 -651 -509 -647
rect -443 -648 -427 -644
rect -110 -642 -90 -636
rect -27 -642 -7 -636
rect 57 -642 77 -636
rect -281 -644 -261 -643
rect -363 -645 -343 -644
rect -359 -649 -343 -645
rect -277 -648 -261 -644
rect -195 -644 -175 -643
rect -191 -648 -175 -644
rect -110 -645 -90 -644
rect -106 -649 -90 -645
rect -27 -645 -7 -644
rect -23 -649 -7 -645
rect 57 -645 77 -644
rect 61 -649 77 -645
rect -608 -658 -592 -654
rect -608 -659 -588 -658
rect -529 -659 -513 -655
rect -447 -656 -431 -652
rect -447 -657 -427 -656
rect -363 -657 -347 -653
rect -281 -656 -265 -652
rect -281 -657 -261 -656
rect -195 -656 -179 -652
rect -195 -657 -175 -656
rect -110 -657 -94 -653
rect -363 -658 -343 -657
rect -529 -660 -509 -659
rect -608 -667 -588 -661
rect -529 -668 -509 -662
rect -447 -665 -427 -659
rect -363 -666 -343 -660
rect -281 -665 -261 -659
rect -110 -658 -90 -657
rect -27 -657 -11 -653
rect -27 -658 -7 -657
rect 57 -657 73 -653
rect 57 -658 77 -657
rect -195 -665 -175 -659
rect -447 -668 -427 -667
rect -608 -670 -588 -669
rect -604 -674 -588 -670
rect -529 -671 -509 -670
rect -525 -675 -509 -671
rect -443 -672 -427 -668
rect -110 -666 -90 -660
rect -27 -666 -7 -660
rect 57 -666 77 -660
rect -281 -668 -261 -667
rect -363 -669 -343 -668
rect -359 -673 -343 -669
rect -277 -672 -261 -668
rect -195 -668 -175 -667
rect -191 -672 -175 -668
rect -110 -669 -90 -668
rect -106 -673 -90 -669
rect -27 -669 -7 -668
rect -23 -673 -7 -669
rect 57 -669 77 -668
rect 61 -673 77 -669
<< ndcontact >>
rect -86 50 -82 54
rect -80 42 -76 46
rect -82 26 -78 30
rect -76 18 -72 22
rect -86 10 -82 14
rect -70 -7 -66 -3
rect -86 -15 -82 -11
rect -70 -32 -66 -28
rect -289 -38 -285 -34
rect -283 -46 -279 -42
rect -82 -42 -78 -38
rect -76 -50 -72 -46
rect -285 -62 -281 -58
rect -279 -70 -275 -66
rect -86 -68 -82 -64
rect -289 -78 -285 -74
rect -70 -76 -66 -72
rect 57 -81 61 -77
rect -273 -95 -269 -91
rect -86 -92 -82 -88
rect 63 -89 67 -85
rect -289 -103 -285 -99
rect -70 -100 -66 -96
rect 61 -105 65 -101
rect 67 -113 71 -109
rect -273 -120 -269 -116
rect 57 -121 61 -117
rect -285 -130 -281 -126
rect -279 -138 -275 -134
rect -41 -139 -37 -135
rect 73 -138 77 -134
rect -35 -147 -31 -143
rect 57 -146 61 -142
rect -491 -158 -487 -154
rect -289 -156 -285 -152
rect -485 -166 -481 -162
rect -273 -164 -269 -160
rect -487 -182 -483 -178
rect -289 -180 -285 -176
rect -481 -190 -477 -186
rect -273 -188 -269 -184
rect -31 -157 -27 -153
rect -37 -166 -33 -162
rect 73 -163 77 -159
rect -31 -175 -27 -171
rect 61 -173 65 -169
rect 67 -181 71 -177
rect -591 -196 -587 -192
rect -491 -198 -487 -194
rect -585 -204 -581 -200
rect -208 -205 -204 -201
rect -147 -189 -143 -185
rect -129 -205 -125 -201
rect -200 -211 -196 -207
rect -475 -215 -471 -211
rect -190 -215 -186 -211
rect -181 -209 -177 -205
rect -172 -215 -168 -211
rect -587 -220 -583 -216
rect -491 -223 -487 -219
rect -392 -220 -388 -216
rect -581 -228 -577 -224
rect -591 -236 -587 -232
rect -398 -228 -394 -224
rect -475 -240 -471 -236
rect -402 -238 -398 -234
rect -575 -253 -571 -249
rect -487 -250 -483 -246
rect -396 -247 -392 -243
rect -591 -261 -587 -257
rect -481 -258 -477 -254
rect -402 -256 -398 -252
rect -575 -278 -571 -274
rect -491 -276 -487 -272
rect -475 -284 -471 -280
rect -587 -288 -583 -284
rect -581 -296 -577 -292
rect -491 -300 -487 -296
rect -475 -308 -471 -304
rect -591 -314 -587 -310
rect -575 -322 -571 -318
rect -304 -286 -300 -282
rect -286 -270 -282 -266
rect 57 -199 61 -195
rect 73 -207 77 -203
rect 57 -223 61 -219
rect 73 -231 77 -227
rect -105 -263 -101 -259
rect -96 -257 -92 -253
rect -54 -259 -50 -255
rect -36 -243 -32 -239
rect -23 -249 -19 -245
rect -15 -243 -11 -239
rect -87 -263 -83 -259
rect -261 -296 -257 -292
rect -252 -290 -248 -286
rect -233 -292 -229 -288
rect -225 -286 -221 -282
rect -243 -296 -239 -292
rect -418 -324 -414 -320
rect -410 -330 -406 -326
rect -397 -324 -393 -320
rect -591 -338 -587 -334
rect 2 -319 6 -315
rect -379 -340 -375 -336
rect -575 -346 -571 -342
rect -346 -344 -342 -340
rect -337 -338 -333 -334
rect -328 -344 -324 -340
rect 10 -325 14 -321
rect 20 -329 24 -325
rect 29 -323 33 -319
rect 38 -329 42 -325
rect -539 -389 -535 -385
rect -531 -383 -527 -379
rect -279 -361 -275 -357
rect -270 -361 -266 -357
rect -262 -367 -258 -363
rect -242 -366 -238 -362
rect -234 -366 -230 -362
rect 54 -339 58 -335
rect 72 -323 76 -319
rect 85 -329 89 -325
rect 93 -323 97 -319
rect 120 -339 124 -335
rect 129 -333 133 -329
rect 148 -335 152 -331
rect 156 -329 160 -325
rect 138 -339 142 -335
rect 179 -351 183 -347
rect 197 -335 201 -331
rect -515 -415 -511 -411
rect -506 -409 -502 -405
rect -487 -411 -483 -407
rect -479 -405 -475 -401
rect -197 -377 -193 -373
rect -189 -383 -185 -379
rect -176 -377 -172 -373
rect 165 -367 169 -363
rect 159 -376 163 -372
rect 165 -385 169 -381
rect -158 -393 -154 -389
rect -497 -415 -493 -411
rect -610 -425 -606 -421
rect -601 -425 -597 -421
rect -593 -431 -589 -427
rect -573 -430 -569 -426
rect -565 -430 -561 -426
rect -466 -427 -462 -423
rect -448 -411 -444 -407
rect -139 -398 -135 -394
rect -130 -392 -126 -388
rect -121 -398 -117 -394
rect -84 -408 -80 -404
rect -76 -408 -72 -404
rect -416 -413 -412 -409
rect -407 -413 -403 -409
rect -399 -419 -395 -415
rect -379 -418 -375 -414
rect -56 -409 -52 -405
rect -48 -403 -44 -399
rect -39 -403 -35 -399
rect -371 -418 -367 -414
rect -564 -462 -560 -458
rect -555 -462 -551 -458
rect -547 -456 -543 -452
rect -500 -452 -496 -448
rect -527 -457 -523 -453
rect -519 -457 -515 -453
rect -491 -458 -487 -454
rect -482 -452 -478 -448
rect -466 -453 -462 -449
rect -404 -462 -400 -458
rect -395 -462 -391 -458
rect -387 -456 -383 -452
rect -340 -452 -336 -448
rect -367 -457 -363 -453
rect -448 -469 -444 -465
rect -359 -457 -355 -453
rect -331 -458 -327 -454
rect -322 -452 -318 -448
rect -306 -453 -302 -449
rect -255 -459 -251 -455
rect -246 -459 -242 -455
rect -238 -453 -234 -449
rect -191 -449 -187 -445
rect -218 -454 -214 -450
rect -288 -469 -284 -465
rect -210 -454 -206 -450
rect -182 -455 -178 -451
rect -173 -449 -169 -445
rect -157 -450 -153 -446
rect -103 -459 -99 -455
rect -94 -459 -90 -455
rect -86 -453 -82 -449
rect -39 -449 -35 -445
rect -66 -454 -62 -450
rect -139 -466 -135 -462
rect -58 -454 -54 -450
rect -30 -455 -26 -451
rect -21 -449 -17 -445
rect -5 -450 -1 -446
rect 13 -466 17 -462
rect 49 -464 53 -460
rect 67 -448 71 -444
rect 83 -464 87 -460
rect 101 -448 105 -444
rect -572 -548 -568 -544
rect -493 -549 -489 -545
rect -411 -546 -407 -542
rect -327 -547 -323 -543
rect -245 -546 -241 -542
rect -159 -546 -155 -542
rect -566 -556 -562 -552
rect -487 -557 -483 -553
rect -74 -547 -70 -543
rect 9 -547 13 -543
rect 93 -547 97 -543
rect -405 -554 -401 -550
rect -321 -555 -317 -551
rect -239 -554 -235 -550
rect -153 -554 -149 -550
rect -68 -555 -64 -551
rect 15 -555 19 -551
rect 99 -555 103 -551
rect -576 -564 -572 -560
rect -497 -565 -493 -561
rect -415 -562 -411 -558
rect -331 -563 -327 -559
rect -249 -562 -245 -558
rect -163 -562 -159 -558
rect -78 -563 -74 -559
rect 5 -563 9 -559
rect 89 -563 93 -559
rect -560 -581 -556 -577
rect -481 -582 -477 -578
rect -399 -579 -395 -575
rect -315 -580 -311 -576
rect -233 -579 -229 -575
rect -147 -579 -143 -575
rect -62 -580 -58 -576
rect 21 -580 25 -576
rect 105 -580 109 -576
rect -576 -589 -572 -585
rect -497 -590 -493 -586
rect -415 -587 -411 -583
rect -331 -588 -327 -584
rect -249 -587 -245 -583
rect -163 -587 -159 -583
rect -78 -588 -74 -584
rect 5 -588 9 -584
rect 89 -588 93 -584
rect -560 -606 -556 -602
rect -481 -607 -477 -603
rect -399 -604 -395 -600
rect -315 -605 -311 -601
rect -233 -604 -229 -600
rect -147 -604 -143 -600
rect -62 -605 -58 -601
rect 21 -605 25 -601
rect 105 -605 109 -601
rect -572 -616 -568 -612
rect -493 -617 -489 -613
rect -411 -614 -407 -610
rect -327 -615 -323 -611
rect -245 -614 -241 -610
rect -159 -614 -155 -610
rect -566 -624 -562 -620
rect -487 -625 -483 -621
rect -74 -615 -70 -611
rect 9 -615 13 -611
rect 93 -615 97 -611
rect -405 -622 -401 -618
rect -321 -623 -317 -619
rect -239 -622 -235 -618
rect -153 -622 -149 -618
rect -68 -623 -64 -619
rect 15 -623 19 -619
rect 99 -623 103 -619
rect -576 -642 -572 -638
rect -497 -643 -493 -639
rect -415 -640 -411 -636
rect -331 -641 -327 -637
rect -249 -640 -245 -636
rect -163 -640 -159 -636
rect -560 -650 -556 -646
rect -481 -651 -477 -647
rect -78 -641 -74 -637
rect 5 -641 9 -637
rect 89 -641 93 -637
rect -399 -648 -395 -644
rect -315 -649 -311 -645
rect -233 -648 -229 -644
rect -147 -648 -143 -644
rect -62 -649 -58 -645
rect 21 -649 25 -645
rect 105 -649 109 -645
rect -576 -666 -572 -662
rect -497 -667 -493 -663
rect -415 -664 -411 -660
rect -331 -665 -327 -661
rect -249 -664 -245 -660
rect -163 -664 -159 -660
rect -560 -674 -556 -670
rect -481 -675 -477 -671
rect -78 -665 -74 -661
rect 5 -665 9 -661
rect 89 -665 93 -661
rect -399 -672 -395 -668
rect -315 -673 -311 -669
rect -233 -672 -229 -668
rect -147 -672 -143 -668
rect -62 -673 -58 -669
rect 21 -673 25 -669
rect 105 -673 109 -669
<< pdcontact >>
rect -102 50 -98 54
rect -118 42 -114 46
rect -102 26 -98 30
rect -118 18 -114 22
rect -102 1 -98 5
rect -118 -7 -114 -3
rect -102 -24 -98 -20
rect -118 -32 -114 -28
rect -305 -38 -301 -34
rect -321 -46 -317 -42
rect -102 -42 -98 -38
rect -118 -50 -114 -46
rect -305 -62 -301 -58
rect -102 -60 -98 -56
rect -321 -70 -317 -66
rect -118 -76 -114 -72
rect -305 -87 -301 -83
rect -102 -84 -98 -80
rect 41 -81 45 -77
rect -321 -95 -317 -91
rect 25 -89 29 -85
rect -118 -100 -114 -96
rect 41 -105 45 -101
rect -305 -112 -301 -108
rect 25 -113 29 -109
rect -321 -120 -317 -116
rect -305 -130 -301 -126
rect 41 -130 45 -126
rect -321 -138 -317 -134
rect -57 -139 -53 -135
rect 25 -138 29 -134
rect -305 -148 -301 -144
rect -73 -147 -69 -143
rect -507 -158 -503 -154
rect -523 -166 -519 -162
rect -321 -164 -317 -160
rect -305 -172 -301 -168
rect -507 -182 -503 -178
rect -523 -190 -519 -186
rect -321 -188 -317 -184
rect -208 -189 -204 -185
rect -200 -173 -196 -169
rect -190 -187 -186 -183
rect -172 -151 -168 -147
rect -147 -151 -143 -147
rect -138 -167 -134 -163
rect -129 -151 -125 -147
rect -59 -157 -55 -153
rect 41 -155 45 -151
rect 25 -163 29 -159
rect -95 -175 -91 -171
rect 41 -173 45 -169
rect 25 -181 29 -177
rect -607 -196 -603 -192
rect -623 -204 -619 -200
rect -507 -207 -503 -203
rect -523 -215 -519 -211
rect 41 -191 45 -187
rect -105 -199 -101 -195
rect -607 -220 -603 -216
rect -376 -220 -372 -216
rect -623 -228 -619 -224
rect -507 -232 -503 -228
rect -360 -228 -356 -224
rect -304 -232 -300 -228
rect -607 -245 -603 -241
rect -523 -240 -519 -236
rect -374 -238 -370 -234
rect -623 -253 -619 -249
rect -507 -250 -503 -246
rect -295 -248 -291 -244
rect -286 -232 -282 -228
rect -261 -232 -257 -228
rect -523 -258 -519 -254
rect -338 -256 -334 -252
rect -607 -270 -603 -266
rect -507 -268 -503 -264
rect -623 -278 -619 -274
rect -523 -284 -519 -280
rect -607 -288 -603 -284
rect -397 -286 -393 -282
rect -623 -296 -619 -292
rect -507 -292 -503 -288
rect -607 -306 -603 -302
rect -523 -308 -519 -304
rect -418 -308 -414 -304
rect -410 -292 -406 -288
rect -388 -302 -384 -298
rect -379 -286 -375 -282
rect -623 -322 -619 -318
rect -346 -316 -342 -312
rect -328 -280 -324 -276
rect -54 -205 -50 -201
rect -45 -221 -41 -217
rect -36 -205 -32 -201
rect 25 -207 29 -203
rect -23 -211 -19 -207
rect -87 -235 -83 -231
rect -243 -268 -239 -264
rect -233 -254 -229 -250
rect 41 -215 45 -211
rect -15 -227 -11 -223
rect 25 -231 29 -227
rect -225 -270 -221 -266
rect 2 -303 6 -299
rect 10 -287 14 -283
rect 20 -301 24 -297
rect 38 -265 42 -261
rect 120 -275 124 -271
rect 54 -285 58 -281
rect 63 -301 67 -297
rect 72 -285 76 -281
rect 85 -291 89 -287
rect -607 -330 -603 -326
rect -623 -346 -619 -342
rect -279 -344 -275 -340
rect -270 -342 -266 -338
rect -262 -328 -258 -324
rect -242 -328 -238 -324
rect 93 -307 97 -303
rect 138 -311 142 -307
rect 148 -297 152 -293
rect -234 -344 -230 -340
rect -176 -339 -172 -335
rect -539 -351 -535 -347
rect -531 -367 -527 -363
rect -515 -351 -511 -347
rect -610 -408 -606 -404
rect -601 -406 -597 -402
rect -593 -392 -589 -388
rect -573 -392 -569 -388
rect -497 -387 -493 -383
rect -487 -373 -483 -369
rect -565 -408 -561 -404
rect -479 -389 -475 -385
rect -466 -373 -462 -369
rect -457 -389 -453 -385
rect -448 -373 -444 -369
rect -197 -361 -193 -357
rect -189 -345 -185 -341
rect -167 -355 -163 -351
rect -158 -339 -154 -335
rect -139 -370 -135 -366
rect -121 -334 -117 -330
rect 156 -313 160 -309
rect 179 -297 183 -293
rect 188 -313 192 -309
rect 197 -297 201 -293
rect -416 -396 -412 -392
rect -407 -394 -403 -390
rect -399 -380 -395 -376
rect -379 -380 -375 -376
rect -371 -396 -367 -392
rect -84 -386 -80 -382
rect -76 -370 -72 -366
rect -56 -370 -52 -366
rect -48 -384 -44 -380
rect 101 -367 105 -363
rect -39 -386 -35 -382
rect 137 -385 141 -381
rect 49 -410 53 -406
rect 58 -426 62 -422
rect 67 -410 71 -406
rect 83 -410 87 -406
rect 92 -426 96 -422
rect 101 -410 105 -406
rect -564 -479 -560 -475
rect -555 -481 -551 -477
rect -547 -495 -543 -491
rect -527 -495 -523 -491
rect -519 -479 -515 -475
rect -500 -516 -496 -512
rect -482 -480 -478 -476
rect -404 -479 -400 -475
rect -466 -507 -462 -503
rect -457 -491 -453 -487
rect -395 -481 -391 -477
rect -387 -495 -383 -491
rect -367 -495 -363 -491
rect -359 -479 -355 -475
rect -448 -507 -444 -503
rect -340 -516 -336 -512
rect -322 -480 -318 -476
rect -255 -476 -251 -472
rect -306 -507 -302 -503
rect -297 -491 -293 -487
rect -246 -478 -242 -474
rect -238 -492 -234 -488
rect -218 -492 -214 -488
rect -210 -476 -206 -472
rect -288 -507 -284 -503
rect -191 -513 -187 -509
rect -173 -477 -169 -473
rect -103 -476 -99 -472
rect -157 -504 -153 -500
rect -148 -488 -144 -484
rect -94 -478 -90 -474
rect -86 -492 -82 -488
rect -66 -492 -62 -488
rect -58 -476 -54 -472
rect -139 -504 -135 -500
rect -39 -513 -35 -509
rect -21 -477 -17 -473
rect -5 -504 -1 -500
rect 4 -488 8 -484
rect 13 -504 17 -500
rect -592 -548 -588 -544
rect -513 -549 -509 -545
rect -431 -546 -427 -542
rect -347 -547 -343 -543
rect -265 -546 -261 -542
rect -179 -546 -175 -542
rect -94 -547 -90 -543
rect -608 -556 -604 -552
rect -529 -557 -525 -553
rect -447 -554 -443 -550
rect -11 -547 -7 -543
rect 73 -547 77 -543
rect -363 -555 -359 -551
rect -281 -554 -277 -550
rect -195 -554 -191 -550
rect -110 -555 -106 -551
rect -27 -555 -23 -551
rect 57 -555 61 -551
rect -592 -573 -588 -569
rect -513 -574 -509 -570
rect -431 -571 -427 -567
rect -347 -572 -343 -568
rect -265 -571 -261 -567
rect -179 -571 -175 -567
rect -94 -572 -90 -568
rect -608 -581 -604 -577
rect -529 -582 -525 -578
rect -447 -579 -443 -575
rect -11 -572 -7 -568
rect 73 -572 77 -568
rect -363 -580 -359 -576
rect -281 -579 -277 -575
rect -195 -579 -191 -575
rect -110 -580 -106 -576
rect -27 -580 -23 -576
rect 57 -580 61 -576
rect -592 -598 -588 -594
rect -513 -599 -509 -595
rect -431 -596 -427 -592
rect -347 -597 -343 -593
rect -265 -596 -261 -592
rect -179 -596 -175 -592
rect -94 -597 -90 -593
rect -608 -606 -604 -602
rect -529 -607 -525 -603
rect -447 -604 -443 -600
rect -11 -597 -7 -593
rect 73 -597 77 -593
rect -363 -605 -359 -601
rect -281 -604 -277 -600
rect -195 -604 -191 -600
rect -110 -605 -106 -601
rect -27 -605 -23 -601
rect 57 -605 61 -601
rect -592 -616 -588 -612
rect -513 -617 -509 -613
rect -431 -614 -427 -610
rect -347 -615 -343 -611
rect -265 -614 -261 -610
rect -179 -614 -175 -610
rect -94 -615 -90 -611
rect -608 -624 -604 -620
rect -529 -625 -525 -621
rect -447 -622 -443 -618
rect -11 -615 -7 -611
rect 73 -615 77 -611
rect -363 -623 -359 -619
rect -281 -622 -277 -618
rect -195 -622 -191 -618
rect -110 -623 -106 -619
rect -27 -623 -23 -619
rect 57 -623 61 -619
rect -592 -634 -588 -630
rect -513 -635 -509 -631
rect -431 -632 -427 -628
rect -347 -633 -343 -629
rect -265 -632 -261 -628
rect -179 -632 -175 -628
rect -94 -633 -90 -629
rect -11 -633 -7 -629
rect 73 -633 77 -629
rect -608 -650 -604 -646
rect -529 -651 -525 -647
rect -447 -648 -443 -644
rect -363 -649 -359 -645
rect -281 -648 -277 -644
rect -195 -648 -191 -644
rect -110 -649 -106 -645
rect -27 -649 -23 -645
rect 57 -649 61 -645
rect -592 -658 -588 -654
rect -513 -659 -509 -655
rect -431 -656 -427 -652
rect -347 -657 -343 -653
rect -265 -656 -261 -652
rect -179 -656 -175 -652
rect -94 -657 -90 -653
rect -11 -657 -7 -653
rect 73 -657 77 -653
rect -608 -674 -604 -670
rect -529 -675 -525 -671
rect -447 -672 -443 -668
rect -363 -673 -359 -669
rect -281 -672 -277 -668
rect -195 -672 -191 -668
rect -110 -673 -106 -669
rect -27 -673 -23 -669
rect 57 -673 61 -669
<< polysilicon >>
rect -122 47 -118 49
rect -98 47 -86 49
rect -76 47 -72 49
rect -122 23 -118 25
rect -98 23 -82 25
rect -72 23 -68 25
rect -90 7 -86 9
rect -66 7 -52 9
rect -121 -2 -118 0
rect -98 -2 -86 0
rect -66 -2 -61 0
rect -90 -18 -86 -16
rect -66 -18 -52 -16
rect -121 -27 -118 -25
rect -98 -27 -86 -25
rect -66 -27 -61 -25
rect -325 -41 -321 -39
rect -301 -41 -289 -39
rect -279 -41 -275 -39
rect -122 -45 -118 -43
rect -98 -45 -82 -43
rect -72 -45 -68 -43
rect -122 -63 -118 -61
rect -98 -63 -54 -61
rect -325 -65 -321 -63
rect -301 -65 -285 -63
rect -275 -65 -271 -63
rect -122 -71 -118 -69
rect -98 -71 -86 -69
rect -66 -71 -63 -69
rect -293 -81 -289 -79
rect -269 -81 -255 -79
rect 21 -84 25 -82
rect 45 -84 57 -82
rect 67 -84 71 -82
rect -122 -87 -118 -85
rect -98 -86 -54 -85
rect -98 -87 -57 -86
rect -324 -90 -321 -88
rect -301 -90 -289 -88
rect -269 -90 -264 -88
rect -122 -95 -118 -93
rect -98 -95 -86 -93
rect -66 -95 -63 -93
rect -293 -106 -289 -104
rect -269 -106 -255 -104
rect 21 -108 25 -106
rect 45 -108 61 -106
rect 71 -108 75 -106
rect -324 -115 -321 -113
rect -301 -115 -289 -113
rect -269 -115 -264 -113
rect 53 -124 57 -122
rect 77 -124 91 -122
rect -325 -133 -321 -131
rect -301 -133 -285 -131
rect -275 -133 -271 -131
rect 22 -133 25 -131
rect 45 -133 57 -131
rect 77 -133 82 -131
rect -76 -142 -73 -140
rect -53 -142 -41 -140
rect -31 -142 -28 -140
rect -185 -147 -183 -144
rect -175 -147 -173 -144
rect -142 -147 -140 -143
rect -132 -147 -130 -143
rect -325 -151 -321 -149
rect -301 -151 -257 -149
rect -325 -159 -321 -157
rect -301 -159 -289 -157
rect -269 -159 -266 -157
rect -527 -161 -523 -159
rect -503 -161 -491 -159
rect -481 -161 -477 -159
rect -203 -169 -201 -166
rect -325 -175 -321 -173
rect -301 -174 -257 -173
rect -301 -175 -260 -174
rect -325 -183 -321 -181
rect -301 -183 -289 -181
rect -269 -183 -266 -181
rect -527 -185 -523 -183
rect -503 -185 -487 -183
rect -477 -185 -473 -183
rect 53 -149 57 -147
rect 77 -149 91 -147
rect 22 -158 25 -156
rect 45 -158 57 -156
rect 77 -158 82 -156
rect -98 -160 -95 -158
rect -55 -160 -37 -158
rect -27 -160 -24 -158
rect -142 -185 -140 -167
rect -132 -185 -130 -167
rect -98 -170 -95 -168
rect -55 -170 -37 -168
rect -27 -170 -24 -168
rect 21 -176 25 -174
rect 45 -176 61 -174
rect 71 -176 75 -174
rect -627 -199 -623 -197
rect -603 -199 -591 -197
rect -581 -199 -577 -197
rect -495 -201 -491 -199
rect -471 -201 -457 -199
rect -203 -201 -201 -189
rect -526 -210 -523 -208
rect -503 -210 -491 -208
rect -471 -210 -466 -208
rect -185 -205 -183 -187
rect -175 -205 -173 -187
rect -100 -195 -98 -192
rect -90 -195 -88 -192
rect 21 -194 25 -192
rect 45 -194 89 -192
rect -203 -214 -201 -211
rect -142 -209 -140 -205
rect -132 -209 -130 -205
rect -627 -223 -623 -221
rect -603 -223 -587 -221
rect -577 -223 -573 -221
rect -185 -218 -183 -215
rect -175 -218 -173 -215
rect -401 -223 -398 -221
rect -388 -223 -376 -221
rect -356 -223 -353 -221
rect -495 -226 -491 -224
rect -471 -226 -457 -224
rect -299 -228 -297 -224
rect -289 -228 -287 -224
rect -256 -228 -254 -225
rect -246 -228 -244 -225
rect -526 -235 -523 -233
rect -503 -235 -491 -233
rect -471 -235 -466 -233
rect -595 -239 -591 -237
rect -571 -239 -557 -237
rect -405 -241 -402 -239
rect -392 -241 -374 -239
rect -334 -241 -331 -239
rect -626 -248 -623 -246
rect -603 -248 -591 -246
rect -571 -248 -566 -246
rect -405 -251 -402 -249
rect -392 -251 -374 -249
rect -334 -251 -331 -249
rect -527 -253 -523 -251
rect -503 -253 -487 -251
rect -477 -253 -473 -251
rect -595 -264 -591 -262
rect -571 -264 -557 -262
rect -299 -266 -297 -248
rect -289 -266 -287 -248
rect -527 -271 -523 -269
rect -503 -271 -459 -269
rect -626 -273 -623 -271
rect -603 -273 -591 -271
rect -571 -273 -566 -271
rect -341 -276 -339 -273
rect -331 -276 -329 -273
rect -527 -279 -523 -277
rect -503 -279 -491 -277
rect -471 -279 -468 -277
rect -392 -282 -390 -278
rect -382 -282 -380 -278
rect -413 -288 -411 -284
rect -627 -291 -623 -289
rect -603 -291 -587 -289
rect -577 -291 -573 -289
rect -527 -295 -523 -293
rect -503 -294 -459 -293
rect -503 -295 -462 -294
rect -527 -303 -523 -301
rect -503 -303 -491 -301
rect -471 -303 -468 -301
rect -627 -309 -623 -307
rect -603 -309 -559 -307
rect -627 -317 -623 -315
rect -603 -317 -591 -315
rect -571 -317 -568 -315
rect -413 -320 -411 -308
rect -392 -320 -390 -302
rect -382 -320 -380 -302
rect -49 -201 -47 -197
rect -39 -201 -37 -197
rect 21 -202 25 -200
rect 45 -202 57 -200
rect 77 -202 80 -200
rect -18 -207 -16 -203
rect -228 -250 -226 -247
rect -256 -286 -254 -268
rect -246 -286 -244 -268
rect -100 -253 -98 -235
rect -90 -253 -88 -235
rect -49 -239 -47 -221
rect -39 -239 -37 -221
rect 21 -218 25 -216
rect 45 -217 89 -216
rect 45 -218 86 -217
rect 21 -226 25 -224
rect 45 -226 57 -224
rect 77 -226 80 -224
rect -18 -239 -16 -227
rect -18 -253 -16 -249
rect -49 -263 -47 -259
rect -39 -263 -37 -259
rect 25 -261 27 -258
rect 35 -261 37 -258
rect -100 -266 -98 -263
rect -90 -266 -88 -263
rect -228 -282 -226 -270
rect -299 -290 -297 -286
rect -289 -290 -287 -286
rect 7 -283 9 -280
rect -228 -295 -226 -292
rect -256 -299 -254 -296
rect -246 -299 -244 -296
rect 125 -271 127 -268
rect 135 -271 137 -268
rect 59 -281 61 -277
rect 69 -281 71 -277
rect 90 -287 92 -283
rect -627 -333 -623 -331
rect -603 -332 -559 -331
rect -603 -333 -562 -332
rect -413 -334 -411 -330
rect -627 -341 -623 -339
rect -603 -341 -591 -339
rect -571 -341 -568 -339
rect -341 -334 -339 -316
rect -331 -334 -329 -316
rect -274 -324 -272 -312
rect 7 -315 9 -303
rect -265 -324 -263 -321
rect -237 -324 -235 -320
rect -534 -347 -532 -343
rect -392 -344 -390 -340
rect -382 -344 -380 -340
rect 25 -319 27 -301
rect 35 -319 37 -301
rect 59 -319 61 -301
rect 69 -319 71 -301
rect 90 -319 92 -307
rect 153 -293 155 -290
rect 184 -293 186 -289
rect 194 -293 196 -289
rect -134 -330 -132 -327
rect -124 -330 -122 -327
rect 7 -328 9 -325
rect -171 -335 -169 -331
rect -161 -335 -159 -331
rect -192 -341 -190 -337
rect -510 -347 -508 -344
rect -500 -347 -498 -344
rect -341 -347 -339 -344
rect -331 -347 -329 -344
rect -605 -388 -603 -376
rect -534 -379 -532 -367
rect -596 -388 -594 -385
rect -568 -388 -566 -384
rect -274 -350 -272 -344
rect -274 -357 -272 -353
rect -265 -357 -263 -344
rect -237 -356 -235 -344
rect -482 -369 -480 -366
rect -461 -369 -459 -365
rect -451 -369 -449 -365
rect -534 -393 -532 -389
rect -510 -405 -508 -387
rect -500 -405 -498 -387
rect -411 -376 -409 -364
rect -274 -369 -272 -367
rect -402 -376 -400 -373
rect -374 -376 -372 -372
rect -274 -373 -273 -369
rect -265 -370 -263 -367
rect -237 -370 -235 -366
rect -192 -373 -190 -361
rect -171 -373 -169 -355
rect -161 -373 -159 -355
rect 25 -332 27 -329
rect 35 -332 37 -329
rect 125 -329 127 -311
rect 135 -329 137 -311
rect 153 -325 155 -313
rect 90 -333 92 -329
rect 184 -331 186 -313
rect 194 -331 196 -313
rect 153 -338 155 -335
rect 59 -343 61 -339
rect 69 -343 71 -339
rect 125 -342 127 -339
rect 135 -342 137 -339
rect -79 -366 -77 -362
rect -51 -366 -49 -363
rect -42 -366 -40 -354
rect 184 -355 186 -351
rect 194 -355 196 -351
rect -274 -374 -272 -373
rect -482 -401 -480 -389
rect -605 -414 -603 -408
rect -605 -421 -603 -417
rect -596 -421 -594 -408
rect -568 -420 -566 -408
rect -461 -407 -459 -389
rect -451 -407 -449 -389
rect -192 -387 -190 -383
rect -134 -388 -132 -370
rect -124 -388 -122 -370
rect 98 -370 101 -368
rect 141 -370 159 -368
rect 169 -370 172 -368
rect 98 -380 101 -378
rect 141 -380 159 -378
rect 169 -380 172 -378
rect -411 -402 -409 -396
rect -482 -414 -480 -411
rect -510 -418 -508 -415
rect -500 -418 -498 -415
rect -411 -409 -409 -405
rect -402 -409 -400 -396
rect -374 -408 -372 -396
rect -171 -397 -169 -393
rect -161 -397 -159 -393
rect -79 -398 -77 -386
rect -134 -401 -132 -398
rect -124 -401 -122 -398
rect -51 -399 -49 -386
rect -42 -392 -40 -386
rect -42 -399 -40 -395
rect -79 -412 -77 -408
rect 54 -406 56 -402
rect 64 -406 66 -402
rect 88 -406 90 -402
rect 98 -406 100 -402
rect -51 -412 -49 -409
rect -42 -411 -40 -409
rect -41 -415 -40 -411
rect -42 -416 -40 -415
rect -411 -421 -409 -419
rect -411 -425 -410 -421
rect -402 -422 -400 -419
rect -374 -422 -372 -418
rect -411 -426 -409 -425
rect -605 -433 -603 -431
rect -605 -437 -604 -433
rect -596 -434 -594 -431
rect -568 -434 -566 -430
rect -461 -431 -459 -427
rect -451 -431 -449 -427
rect -605 -438 -603 -437
rect -250 -443 -248 -442
rect -559 -446 -557 -445
rect -559 -450 -558 -446
rect -495 -448 -493 -445
rect -485 -448 -483 -445
rect -559 -452 -557 -450
rect -550 -452 -548 -449
rect -522 -453 -520 -449
rect -559 -466 -557 -462
rect -559 -475 -557 -469
rect -550 -475 -548 -462
rect -461 -449 -459 -445
rect -451 -449 -449 -445
rect -399 -446 -397 -445
rect -522 -475 -520 -463
rect -495 -476 -493 -458
rect -485 -476 -483 -458
rect -399 -450 -398 -446
rect -335 -448 -333 -445
rect -325 -448 -323 -445
rect -399 -452 -397 -450
rect -390 -452 -388 -449
rect -362 -453 -360 -449
rect -399 -466 -397 -462
rect -559 -507 -557 -495
rect -550 -498 -548 -495
rect -522 -499 -520 -495
rect -461 -487 -459 -469
rect -451 -487 -449 -469
rect -399 -475 -397 -469
rect -390 -475 -388 -462
rect -301 -449 -299 -445
rect -291 -449 -289 -445
rect -250 -447 -249 -443
rect -186 -445 -184 -442
rect -176 -445 -174 -442
rect -250 -449 -248 -447
rect -241 -449 -239 -446
rect -362 -475 -360 -463
rect -335 -476 -333 -458
rect -325 -476 -323 -458
rect -213 -450 -211 -446
rect -250 -463 -248 -459
rect -399 -507 -397 -495
rect -390 -498 -388 -495
rect -362 -499 -360 -495
rect -461 -511 -459 -507
rect -451 -511 -449 -507
rect -301 -487 -299 -469
rect -291 -487 -289 -469
rect -250 -472 -248 -466
rect -241 -472 -239 -459
rect -152 -446 -150 -442
rect -142 -446 -140 -442
rect -98 -443 -96 -442
rect -213 -472 -211 -460
rect -186 -473 -184 -455
rect -176 -473 -174 -455
rect -98 -447 -97 -443
rect -34 -445 -32 -442
rect -24 -445 -22 -442
rect -98 -449 -96 -447
rect -89 -449 -87 -446
rect -61 -450 -59 -446
rect -98 -463 -96 -459
rect -250 -504 -248 -492
rect -241 -495 -239 -492
rect -213 -496 -211 -492
rect -301 -511 -299 -507
rect -291 -511 -289 -507
rect -152 -484 -150 -466
rect -142 -484 -140 -466
rect -98 -472 -96 -466
rect -89 -472 -87 -459
rect 0 -446 2 -442
rect 10 -446 12 -442
rect 54 -444 56 -426
rect 64 -444 66 -426
rect 88 -444 90 -426
rect 98 -444 100 -426
rect -61 -472 -59 -460
rect -34 -473 -32 -455
rect -24 -473 -22 -455
rect -98 -504 -96 -492
rect -89 -495 -87 -492
rect -61 -496 -59 -492
rect -152 -508 -150 -504
rect -142 -508 -140 -504
rect 0 -484 2 -466
rect 10 -484 12 -466
rect 54 -468 56 -464
rect 64 -468 66 -464
rect 88 -468 90 -464
rect 98 -468 100 -464
rect 0 -508 2 -504
rect 10 -508 12 -504
rect -186 -516 -184 -513
rect -176 -516 -174 -513
rect -34 -516 -32 -513
rect -24 -516 -22 -513
rect -495 -519 -493 -516
rect -485 -519 -483 -516
rect -335 -519 -333 -516
rect -325 -519 -323 -516
rect -612 -551 -608 -549
rect -588 -551 -572 -549
rect -562 -551 -558 -549
rect -451 -549 -447 -547
rect -427 -549 -411 -547
rect -401 -549 -397 -547
rect -533 -552 -529 -550
rect -509 -552 -493 -550
rect -483 -552 -479 -550
rect -367 -550 -363 -548
rect -343 -550 -327 -548
rect -317 -550 -313 -548
rect -285 -549 -281 -547
rect -261 -549 -245 -547
rect -235 -549 -231 -547
rect -199 -549 -195 -547
rect -175 -549 -159 -547
rect -149 -549 -145 -547
rect -114 -550 -110 -548
rect -90 -550 -74 -548
rect -64 -550 -60 -548
rect -31 -550 -27 -548
rect -7 -550 9 -548
rect 19 -550 23 -548
rect 53 -550 57 -548
rect 77 -550 93 -548
rect 103 -550 107 -548
rect -419 -565 -415 -563
rect -395 -565 -381 -563
rect -580 -567 -576 -565
rect -556 -567 -542 -565
rect -501 -568 -497 -566
rect -477 -568 -463 -566
rect -611 -576 -608 -574
rect -588 -576 -576 -574
rect -556 -576 -551 -574
rect -335 -566 -331 -564
rect -311 -566 -297 -564
rect -253 -565 -249 -563
rect -229 -565 -215 -563
rect -167 -565 -163 -563
rect -143 -565 -129 -563
rect -450 -574 -447 -572
rect -427 -574 -415 -572
rect -395 -574 -390 -572
rect -82 -566 -78 -564
rect -58 -566 -44 -564
rect 1 -566 5 -564
rect 25 -566 39 -564
rect 85 -566 89 -564
rect 109 -566 123 -564
rect -532 -577 -529 -575
rect -509 -577 -497 -575
rect -477 -577 -472 -575
rect -366 -575 -363 -573
rect -343 -575 -331 -573
rect -311 -575 -306 -573
rect -284 -574 -281 -572
rect -261 -574 -249 -572
rect -229 -574 -224 -572
rect -198 -574 -195 -572
rect -175 -574 -163 -572
rect -143 -574 -138 -572
rect -113 -575 -110 -573
rect -90 -575 -78 -573
rect -58 -575 -53 -573
rect -30 -575 -27 -573
rect -7 -575 5 -573
rect 25 -575 30 -573
rect 54 -575 57 -573
rect 77 -575 89 -573
rect 109 -575 114 -573
rect -419 -590 -415 -588
rect -395 -590 -381 -588
rect -580 -592 -576 -590
rect -556 -592 -542 -590
rect -501 -593 -497 -591
rect -477 -593 -463 -591
rect -611 -601 -608 -599
rect -588 -601 -576 -599
rect -556 -601 -551 -599
rect -335 -591 -331 -589
rect -311 -591 -297 -589
rect -253 -590 -249 -588
rect -229 -590 -215 -588
rect -167 -590 -163 -588
rect -143 -590 -129 -588
rect -450 -599 -447 -597
rect -427 -599 -415 -597
rect -395 -599 -390 -597
rect -82 -591 -78 -589
rect -58 -591 -44 -589
rect 1 -591 5 -589
rect 25 -591 39 -589
rect 85 -591 89 -589
rect 109 -591 123 -589
rect -532 -602 -529 -600
rect -509 -602 -497 -600
rect -477 -602 -472 -600
rect -366 -600 -363 -598
rect -343 -600 -331 -598
rect -311 -600 -306 -598
rect -284 -599 -281 -597
rect -261 -599 -249 -597
rect -229 -599 -224 -597
rect -198 -599 -195 -597
rect -175 -599 -163 -597
rect -143 -599 -138 -597
rect -113 -600 -110 -598
rect -90 -600 -78 -598
rect -58 -600 -53 -598
rect -30 -600 -27 -598
rect -7 -600 5 -598
rect 25 -600 30 -598
rect 54 -600 57 -598
rect 77 -600 89 -598
rect 109 -600 114 -598
rect -612 -619 -608 -617
rect -588 -619 -572 -617
rect -562 -619 -558 -617
rect -451 -617 -447 -615
rect -427 -617 -411 -615
rect -401 -617 -397 -615
rect -533 -620 -529 -618
rect -509 -620 -493 -618
rect -483 -620 -479 -618
rect -367 -618 -363 -616
rect -343 -618 -327 -616
rect -317 -618 -313 -616
rect -285 -617 -281 -615
rect -261 -617 -245 -615
rect -235 -617 -231 -615
rect -199 -617 -195 -615
rect -175 -617 -159 -615
rect -149 -617 -145 -615
rect -114 -618 -110 -616
rect -90 -618 -74 -616
rect -64 -618 -60 -616
rect -31 -618 -27 -616
rect -7 -618 9 -616
rect 19 -618 23 -616
rect 53 -618 57 -616
rect 77 -618 93 -616
rect 103 -618 107 -616
rect -451 -635 -447 -633
rect -427 -635 -383 -633
rect -612 -637 -608 -635
rect -588 -637 -544 -635
rect -533 -638 -529 -636
rect -509 -638 -465 -636
rect -612 -645 -608 -643
rect -588 -645 -576 -643
rect -556 -645 -553 -643
rect -367 -636 -363 -634
rect -343 -636 -299 -634
rect -285 -635 -281 -633
rect -261 -635 -217 -633
rect -199 -635 -195 -633
rect -175 -635 -131 -633
rect -451 -643 -447 -641
rect -427 -643 -415 -641
rect -395 -643 -392 -641
rect -114 -636 -110 -634
rect -90 -636 -46 -634
rect -31 -636 -27 -634
rect -7 -636 37 -634
rect 53 -636 57 -634
rect 77 -636 121 -634
rect -533 -646 -529 -644
rect -509 -646 -497 -644
rect -477 -646 -474 -644
rect -367 -644 -363 -642
rect -343 -644 -331 -642
rect -311 -644 -308 -642
rect -285 -643 -281 -641
rect -261 -643 -249 -641
rect -229 -643 -226 -641
rect -199 -643 -195 -641
rect -175 -643 -163 -641
rect -143 -643 -140 -641
rect -114 -644 -110 -642
rect -90 -644 -78 -642
rect -58 -644 -55 -642
rect -31 -644 -27 -642
rect -7 -644 5 -642
rect 25 -644 28 -642
rect 53 -644 57 -642
rect 77 -644 89 -642
rect 109 -644 112 -642
rect -451 -659 -447 -657
rect -427 -658 -383 -657
rect -427 -659 -386 -658
rect -612 -661 -608 -659
rect -588 -660 -544 -659
rect -588 -661 -547 -660
rect -533 -662 -529 -660
rect -509 -661 -465 -660
rect -509 -662 -468 -661
rect -612 -669 -608 -667
rect -588 -669 -576 -667
rect -556 -669 -553 -667
rect -367 -660 -363 -658
rect -343 -659 -299 -658
rect -285 -659 -281 -657
rect -261 -658 -217 -657
rect -261 -659 -220 -658
rect -343 -660 -302 -659
rect -451 -667 -447 -665
rect -427 -667 -415 -665
rect -395 -667 -392 -665
rect -199 -659 -195 -657
rect -175 -658 -131 -657
rect -175 -659 -134 -658
rect -114 -660 -110 -658
rect -90 -659 -46 -658
rect -90 -660 -49 -659
rect -533 -670 -529 -668
rect -509 -670 -497 -668
rect -477 -670 -474 -668
rect -367 -668 -363 -666
rect -343 -668 -331 -666
rect -311 -668 -308 -666
rect -285 -667 -281 -665
rect -261 -667 -249 -665
rect -229 -667 -226 -665
rect -199 -667 -195 -665
rect -175 -667 -163 -665
rect -143 -667 -140 -665
rect -31 -660 -27 -658
rect -7 -659 37 -658
rect -7 -660 34 -659
rect 53 -660 57 -658
rect 77 -659 121 -658
rect 77 -660 118 -659
rect -114 -668 -110 -666
rect -90 -668 -78 -666
rect -58 -668 -55 -666
rect -31 -668 -27 -666
rect -7 -668 5 -666
rect 25 -668 28 -666
rect 53 -668 57 -666
rect 77 -668 89 -666
rect 109 -668 112 -666
<< polycontact >>
rect -91 43 -87 47
rect -90 19 -86 23
rect -57 3 -53 7
rect -91 -6 -87 -2
rect -57 -22 -53 -18
rect -91 -31 -87 -27
rect -294 -45 -290 -41
rect -90 -49 -86 -45
rect -293 -69 -289 -65
rect -57 -67 -53 -63
rect -91 -75 -87 -71
rect -260 -85 -256 -81
rect -294 -94 -290 -90
rect -57 -90 -53 -86
rect 52 -88 56 -84
rect -91 -99 -87 -95
rect -260 -110 -256 -106
rect 53 -112 57 -108
rect -294 -119 -290 -115
rect 86 -128 90 -124
rect -293 -137 -289 -133
rect 52 -137 56 -133
rect -46 -146 -42 -142
rect -260 -155 -256 -151
rect -496 -165 -492 -161
rect -294 -163 -290 -159
rect -260 -178 -256 -174
rect -495 -189 -491 -185
rect -294 -187 -290 -183
rect 86 -153 90 -149
rect -140 -184 -136 -180
rect -48 -164 -44 -160
rect 52 -162 56 -158
rect -130 -178 -126 -174
rect -42 -174 -38 -170
rect 53 -180 57 -176
rect -596 -203 -592 -199
rect -201 -200 -197 -196
rect -462 -205 -458 -201
rect -496 -214 -492 -210
rect -183 -198 -179 -194
rect -173 -204 -169 -200
rect -595 -227 -591 -223
rect -462 -230 -458 -226
rect -387 -227 -383 -223
rect -562 -243 -558 -239
rect -496 -239 -492 -235
rect -596 -252 -592 -248
rect -385 -245 -381 -241
rect -495 -257 -491 -253
rect -391 -255 -387 -251
rect -303 -259 -299 -255
rect -562 -268 -558 -264
rect -293 -265 -289 -261
rect -596 -277 -592 -273
rect -462 -275 -458 -271
rect -496 -283 -492 -279
rect -595 -295 -591 -291
rect -462 -298 -458 -294
rect -496 -307 -492 -303
rect -562 -313 -558 -309
rect -596 -321 -592 -317
rect -411 -319 -407 -315
rect -390 -319 -386 -315
rect -380 -313 -376 -309
rect 86 -198 90 -194
rect 52 -206 56 -202
rect -53 -232 -49 -228
rect -260 -285 -256 -281
rect -250 -279 -246 -275
rect -104 -252 -100 -248
rect -94 -246 -90 -242
rect -43 -238 -39 -234
rect 86 -221 90 -217
rect -22 -238 -18 -234
rect 52 -230 56 -226
rect -232 -281 -228 -277
rect -562 -336 -558 -332
rect -339 -327 -335 -323
rect -272 -317 -268 -313
rect 9 -314 13 -310
rect -329 -333 -325 -329
rect -596 -345 -592 -341
rect 27 -312 31 -308
rect 55 -311 59 -307
rect 37 -318 41 -314
rect 65 -318 69 -314
rect 86 -318 90 -314
rect -603 -381 -599 -377
rect -538 -378 -534 -374
rect -263 -355 -259 -351
rect -241 -355 -237 -351
rect -514 -404 -510 -400
rect -504 -398 -500 -394
rect -409 -369 -405 -365
rect -273 -373 -269 -369
rect -190 -372 -186 -368
rect -169 -372 -165 -368
rect -159 -366 -155 -362
rect 121 -328 125 -324
rect 131 -322 135 -318
rect 149 -324 153 -320
rect 180 -324 184 -320
rect 190 -330 194 -326
rect -46 -359 -42 -355
rect -486 -400 -482 -396
rect -465 -400 -461 -396
rect -594 -419 -590 -415
rect -572 -419 -568 -415
rect -455 -406 -451 -402
rect -132 -381 -128 -377
rect -122 -387 -118 -383
rect 154 -368 158 -364
rect 148 -378 152 -374
rect -400 -407 -396 -403
rect -378 -407 -374 -403
rect -77 -397 -73 -393
rect -55 -397 -51 -393
rect -45 -415 -41 -411
rect -410 -425 -406 -421
rect -604 -437 -600 -433
rect 50 -437 54 -433
rect -558 -450 -554 -446
rect -499 -463 -495 -459
rect -548 -468 -544 -464
rect -526 -468 -522 -464
rect -489 -469 -485 -465
rect -398 -450 -394 -446
rect -557 -506 -553 -502
rect -465 -480 -461 -476
rect -455 -474 -451 -470
rect -249 -447 -245 -443
rect -339 -463 -335 -459
rect -388 -468 -384 -464
rect -366 -468 -362 -464
rect -329 -469 -325 -465
rect -397 -506 -393 -502
rect -305 -480 -301 -476
rect -295 -474 -291 -470
rect -190 -460 -186 -456
rect -239 -465 -235 -461
rect -217 -465 -213 -461
rect -180 -466 -176 -462
rect -97 -447 -93 -443
rect -248 -503 -244 -499
rect -156 -477 -152 -473
rect -146 -471 -142 -467
rect 60 -443 64 -439
rect 84 -437 88 -433
rect 94 -443 98 -439
rect -38 -460 -34 -456
rect -87 -465 -83 -461
rect -65 -465 -61 -461
rect -28 -466 -24 -462
rect -96 -503 -92 -499
rect -4 -477 0 -473
rect 6 -471 10 -467
rect -580 -555 -576 -551
rect -501 -556 -497 -552
rect -419 -553 -415 -549
rect -335 -554 -331 -550
rect -253 -553 -249 -549
rect -167 -553 -163 -549
rect -82 -554 -78 -550
rect 1 -554 5 -550
rect 85 -554 89 -550
rect -547 -571 -543 -567
rect -468 -572 -464 -568
rect -386 -569 -382 -565
rect -302 -570 -298 -566
rect -220 -569 -216 -565
rect -134 -569 -130 -565
rect -581 -580 -577 -576
rect -502 -581 -498 -577
rect -420 -578 -416 -574
rect -49 -570 -45 -566
rect 34 -570 38 -566
rect 118 -570 122 -566
rect -336 -579 -332 -575
rect -254 -578 -250 -574
rect -168 -578 -164 -574
rect -83 -579 -79 -575
rect 0 -579 4 -575
rect 84 -579 88 -575
rect -547 -596 -543 -592
rect -468 -597 -464 -593
rect -386 -594 -382 -590
rect -302 -595 -298 -591
rect -220 -594 -216 -590
rect -134 -594 -130 -590
rect -581 -605 -577 -601
rect -502 -606 -498 -602
rect -420 -603 -416 -599
rect -49 -595 -45 -591
rect 34 -595 38 -591
rect 118 -595 122 -591
rect -336 -604 -332 -600
rect -254 -603 -250 -599
rect -168 -603 -164 -599
rect -83 -604 -79 -600
rect 0 -604 4 -600
rect 84 -604 88 -600
rect -580 -623 -576 -619
rect -501 -624 -497 -620
rect -419 -621 -415 -617
rect -335 -622 -331 -618
rect -253 -621 -249 -617
rect -167 -621 -163 -617
rect -82 -622 -78 -618
rect 1 -622 5 -618
rect 85 -622 89 -618
rect -547 -641 -543 -637
rect -468 -642 -464 -638
rect -386 -639 -382 -635
rect -302 -640 -298 -636
rect -220 -639 -216 -635
rect -134 -639 -130 -635
rect -581 -649 -577 -645
rect -502 -650 -498 -646
rect -420 -647 -416 -643
rect -49 -640 -45 -636
rect 34 -640 38 -636
rect 118 -640 122 -636
rect -336 -648 -332 -644
rect -254 -647 -250 -643
rect -168 -647 -164 -643
rect -83 -648 -79 -644
rect 0 -648 4 -644
rect 84 -648 88 -644
rect -547 -664 -543 -660
rect -468 -665 -464 -661
rect -386 -662 -382 -658
rect -302 -663 -298 -659
rect -220 -662 -216 -658
rect -134 -662 -130 -658
rect -581 -673 -577 -669
rect -502 -674 -498 -670
rect -420 -671 -416 -667
rect -49 -663 -45 -659
rect 34 -663 38 -659
rect 118 -663 122 -659
rect -336 -672 -332 -668
rect -254 -671 -250 -667
rect -168 -671 -164 -667
rect -83 -672 -79 -668
rect 0 -672 4 -668
rect 84 -672 88 -668
<< metal1 >>
rect -128 45 -125 61
rect -91 54 -88 58
rect -98 51 -86 54
rect -128 42 -118 45
rect -128 21 -125 42
rect -91 33 -88 43
rect -71 45 -68 61
rect -76 42 -68 45
rect -71 36 -68 42
rect -91 30 -87 33
rect -98 26 -82 30
rect -128 18 -118 21
rect -128 -4 -125 18
rect -90 14 -87 19
rect -72 18 -60 21
rect -101 11 -86 14
rect -101 5 -98 11
rect -128 -7 -118 -4
rect -331 -43 -328 -27
rect -294 -34 -291 -30
rect -301 -37 -289 -34
rect -331 -46 -321 -43
rect -331 -67 -328 -46
rect -294 -55 -291 -45
rect -274 -43 -271 -27
rect -279 -46 -271 -43
rect -274 -52 -271 -46
rect -128 -29 -125 -7
rect -90 -11 -87 -6
rect -63 -4 -60 18
rect -66 -7 -60 -4
rect -101 -14 -86 -11
rect -101 -20 -98 -14
rect -128 -32 -118 -29
rect -128 -47 -125 -32
rect -90 -38 -87 -31
rect -63 -29 -60 -7
rect -56 -18 -53 3
rect -66 -32 -60 -29
rect -98 -42 -82 -38
rect -128 -50 -118 -47
rect -294 -58 -290 -55
rect -301 -62 -285 -58
rect -331 -70 -321 -67
rect -331 -92 -328 -70
rect -293 -74 -290 -69
rect -275 -70 -263 -67
rect -304 -77 -289 -74
rect -304 -83 -301 -77
rect -331 -95 -321 -92
rect -331 -117 -328 -95
rect -293 -99 -290 -94
rect -266 -92 -263 -70
rect -128 -73 -125 -50
rect -90 -56 -87 -49
rect -63 -47 -60 -32
rect -72 -50 -60 -47
rect -98 -59 -87 -56
rect -90 -64 -87 -59
rect -90 -67 -86 -64
rect -128 -76 -118 -73
rect -269 -95 -263 -92
rect -304 -102 -289 -99
rect -304 -108 -301 -102
rect -331 -120 -321 -117
rect -331 -135 -328 -120
rect -293 -126 -290 -119
rect -266 -117 -263 -95
rect -259 -106 -256 -85
rect -128 -97 -125 -76
rect -90 -80 -87 -75
rect -63 -73 -60 -50
rect -56 -63 -53 -22
rect -66 -76 -60 -73
rect -98 -83 -87 -80
rect -90 -88 -87 -83
rect -90 -91 -86 -88
rect -128 -100 -118 -97
rect -90 -103 -87 -99
rect -63 -97 -60 -76
rect -56 -86 -53 -67
rect -66 -100 -60 -97
rect -56 -106 -53 -90
rect 15 -86 18 -70
rect 52 -77 55 -73
rect 45 -80 57 -77
rect 15 -89 25 -86
rect -269 -120 -263 -117
rect -301 -130 -285 -126
rect -331 -138 -321 -135
rect -533 -163 -530 -147
rect -496 -154 -493 -150
rect -503 -157 -491 -154
rect -533 -166 -523 -163
rect -633 -201 -630 -185
rect -596 -192 -593 -188
rect -603 -195 -591 -192
rect -633 -204 -623 -201
rect -633 -225 -630 -204
rect -596 -213 -593 -203
rect -576 -201 -573 -185
rect -581 -204 -573 -201
rect -576 -210 -573 -204
rect -533 -187 -530 -166
rect -496 -175 -493 -165
rect -476 -163 -473 -147
rect -481 -166 -473 -163
rect -476 -172 -473 -166
rect -331 -161 -328 -138
rect -293 -144 -290 -137
rect -266 -135 -263 -120
rect -275 -138 -263 -135
rect -301 -147 -290 -144
rect -293 -152 -290 -147
rect -293 -155 -289 -152
rect -331 -164 -321 -161
rect -496 -178 -492 -175
rect -503 -182 -487 -178
rect -331 -185 -328 -164
rect -293 -168 -290 -163
rect -266 -161 -263 -138
rect -259 -151 -256 -110
rect 15 -110 18 -89
rect 52 -98 55 -88
rect 72 -86 75 -70
rect 67 -89 75 -86
rect 72 -95 75 -89
rect 52 -101 56 -98
rect 45 -105 61 -101
rect 15 -113 25 -110
rect -83 -131 -43 -128
rect -269 -164 -263 -161
rect -301 -171 -290 -168
rect -293 -176 -290 -171
rect -293 -179 -289 -176
rect -533 -190 -523 -187
rect -533 -212 -530 -190
rect -495 -194 -492 -189
rect -477 -190 -465 -187
rect -331 -188 -321 -185
rect -506 -197 -491 -194
rect -506 -203 -503 -197
rect -596 -216 -592 -213
rect -533 -215 -523 -212
rect -603 -220 -587 -216
rect -633 -228 -623 -225
rect -633 -250 -630 -228
rect -595 -232 -592 -227
rect -577 -228 -565 -225
rect -606 -235 -591 -232
rect -606 -241 -603 -235
rect -633 -253 -623 -250
rect -633 -275 -630 -253
rect -595 -257 -592 -252
rect -568 -250 -565 -228
rect -533 -237 -530 -215
rect -495 -219 -492 -214
rect -468 -212 -465 -190
rect -293 -191 -290 -187
rect -266 -185 -263 -164
rect -259 -174 -256 -155
rect -199 -140 -124 -137
rect -83 -137 -80 -131
rect -46 -135 -43 -131
rect 15 -135 18 -113
rect 53 -117 56 -112
rect 71 -113 83 -110
rect 42 -120 57 -117
rect 42 -126 45 -120
rect -111 -140 -80 -137
rect -53 -138 -41 -135
rect 15 -138 25 -135
rect -199 -158 -196 -140
rect -171 -147 -168 -140
rect -147 -147 -143 -140
rect -128 -147 -125 -140
rect -269 -188 -263 -185
rect -259 -194 -256 -178
rect -223 -161 -196 -158
rect -471 -215 -465 -212
rect -506 -222 -491 -219
rect -506 -228 -503 -222
rect -571 -253 -565 -250
rect -606 -260 -591 -257
rect -606 -266 -603 -260
rect -633 -278 -623 -275
rect -633 -293 -630 -278
rect -595 -284 -592 -277
rect -568 -275 -565 -253
rect -561 -264 -558 -243
rect -571 -278 -565 -275
rect -603 -288 -587 -284
rect -633 -296 -623 -293
rect -633 -319 -630 -296
rect -595 -302 -592 -295
rect -568 -293 -565 -278
rect -577 -296 -565 -293
rect -603 -305 -592 -302
rect -595 -310 -592 -305
rect -595 -313 -591 -310
rect -633 -322 -623 -319
rect -633 -343 -630 -322
rect -595 -326 -592 -321
rect -568 -319 -565 -296
rect -561 -309 -558 -268
rect -533 -240 -523 -237
rect -533 -255 -530 -240
rect -495 -246 -492 -239
rect -468 -237 -465 -215
rect -461 -226 -458 -205
rect -386 -212 -346 -209
rect -386 -216 -383 -212
rect -388 -219 -376 -216
rect -349 -218 -346 -212
rect -349 -221 -318 -218
rect -223 -218 -220 -161
rect -199 -169 -196 -161
rect -138 -168 -135 -167
rect -147 -171 -135 -168
rect -147 -180 -144 -171
rect -111 -174 -108 -140
rect -126 -177 -108 -174
rect -100 -147 -73 -144
rect -105 -172 -102 -149
rect -46 -153 -43 -146
rect -31 -147 -20 -144
rect -23 -153 -20 -147
rect -55 -156 -38 -153
rect -41 -162 -38 -156
rect -27 -156 -20 -153
rect -105 -175 -95 -172
rect -165 -183 -144 -180
rect -208 -196 -205 -189
rect -190 -196 -187 -187
rect -165 -194 -162 -183
rect -147 -185 -144 -183
rect -136 -184 -117 -181
rect -120 -187 -117 -184
rect -105 -185 -102 -175
rect -48 -181 -45 -164
rect -41 -165 -37 -162
rect -23 -171 -20 -156
rect 15 -160 18 -138
rect 53 -142 56 -137
rect 80 -135 83 -113
rect 77 -138 83 -135
rect 42 -145 57 -142
rect 42 -151 45 -145
rect 15 -163 25 -160
rect -42 -176 -38 -174
rect -27 -175 -23 -172
rect -42 -178 -41 -176
rect 15 -178 18 -163
rect 53 -169 56 -162
rect 80 -160 83 -138
rect 87 -149 90 -128
rect 77 -163 83 -160
rect 45 -173 61 -169
rect 15 -181 25 -178
rect -105 -188 -57 -185
rect -210 -201 -205 -196
rect -197 -199 -187 -196
rect -179 -197 -162 -194
rect -105 -195 -102 -188
rect -60 -191 -57 -188
rect -60 -194 4 -191
rect -190 -201 -187 -199
rect -190 -204 -178 -201
rect -169 -203 -165 -200
rect -181 -205 -178 -204
rect -54 -201 -51 -194
rect -36 -201 -32 -194
rect -128 -210 -125 -205
rect -23 -207 -20 -194
rect -305 -221 -220 -218
rect -199 -219 -196 -211
rect -190 -219 -187 -215
rect -171 -219 -168 -215
rect -164 -213 -116 -210
rect -164 -219 -161 -213
rect -471 -240 -465 -237
rect -503 -250 -487 -246
rect -533 -258 -523 -255
rect -533 -281 -530 -258
rect -495 -264 -492 -257
rect -468 -255 -465 -240
rect -477 -258 -465 -255
rect -503 -267 -492 -264
rect -495 -272 -492 -267
rect -495 -275 -491 -272
rect -533 -284 -523 -281
rect -533 -305 -530 -284
rect -495 -288 -492 -283
rect -468 -281 -465 -258
rect -461 -271 -458 -230
rect -409 -228 -398 -225
rect -409 -234 -406 -228
rect -386 -234 -383 -227
rect -356 -228 -329 -225
rect -409 -237 -402 -234
rect -409 -252 -406 -237
rect -391 -237 -374 -234
rect -391 -243 -388 -237
rect -392 -246 -388 -243
rect -406 -256 -402 -253
rect -390 -260 -387 -255
rect -438 -264 -387 -260
rect -384 -262 -381 -245
rect -327 -253 -324 -230
rect -334 -256 -324 -253
rect -327 -266 -324 -256
rect -321 -255 -318 -221
rect -304 -228 -301 -221
rect -286 -228 -282 -221
rect -261 -228 -258 -221
rect -294 -249 -291 -248
rect -294 -252 -282 -249
rect -321 -258 -303 -255
rect -285 -261 -282 -252
rect -233 -250 -230 -221
rect -208 -222 -161 -219
rect -372 -269 -324 -266
rect -307 -265 -293 -262
rect -285 -264 -264 -261
rect -285 -266 -282 -264
rect -372 -272 -369 -269
rect -471 -284 -465 -281
rect -503 -291 -492 -288
rect -495 -296 -492 -291
rect -495 -299 -491 -296
rect -533 -308 -523 -305
rect -495 -311 -492 -307
rect -468 -305 -465 -284
rect -461 -294 -458 -275
rect -471 -308 -465 -305
rect -571 -322 -565 -319
rect -603 -329 -592 -326
rect -595 -334 -592 -329
rect -595 -337 -591 -334
rect -633 -346 -623 -343
rect -595 -349 -592 -345
rect -568 -343 -565 -322
rect -561 -332 -558 -313
rect -461 -314 -458 -298
rect -448 -275 -369 -272
rect -571 -346 -565 -343
rect -561 -352 -558 -336
rect -555 -338 -484 -337
rect -555 -340 -472 -338
rect -555 -341 -545 -340
rect -555 -368 -551 -341
rect -539 -347 -536 -340
rect -515 -347 -512 -340
rect -487 -341 -472 -340
rect -487 -359 -484 -341
rect -475 -348 -472 -341
rect -448 -348 -445 -275
rect -409 -288 -406 -275
rect -397 -282 -393 -275
rect -378 -282 -375 -275
rect -327 -276 -324 -269
rect -267 -275 -264 -264
rect -267 -278 -250 -275
rect -242 -277 -239 -268
rect -224 -277 -221 -270
rect -242 -280 -232 -277
rect -264 -284 -260 -281
rect -242 -282 -239 -280
rect -224 -280 -218 -277
rect -224 -282 -221 -280
rect -251 -285 -239 -282
rect -251 -286 -248 -285
rect -304 -291 -301 -286
rect -313 -294 -265 -291
rect -388 -303 -385 -302
rect -397 -306 -385 -303
rect -418 -315 -415 -308
rect -397 -315 -394 -306
rect -376 -312 -349 -309
rect -421 -318 -415 -315
rect -418 -320 -415 -318
rect -407 -318 -394 -315
rect -397 -320 -394 -318
rect -386 -319 -372 -316
rect -352 -325 -349 -312
rect -346 -325 -343 -316
rect -352 -328 -343 -325
rect -335 -326 -322 -323
rect -409 -344 -406 -330
rect -346 -330 -343 -328
rect -346 -333 -334 -330
rect -325 -332 -317 -329
rect -337 -334 -334 -333
rect -412 -347 -410 -344
rect -475 -351 -445 -348
rect -378 -345 -375 -340
rect -405 -348 -369 -345
rect -346 -348 -343 -344
rect -327 -348 -324 -344
rect -313 -348 -310 -294
rect -268 -300 -265 -294
rect -261 -300 -258 -296
rect -242 -300 -239 -296
rect -233 -300 -230 -292
rect -208 -300 -205 -222
rect -119 -267 -116 -213
rect -44 -222 -41 -221
rect -44 -225 -32 -222
rect -80 -231 -53 -228
rect -107 -245 -94 -242
rect -86 -244 -83 -235
rect -80 -244 -77 -231
rect -35 -234 -32 -225
rect -14 -234 -11 -227
rect -67 -238 -43 -235
rect -35 -237 -22 -234
rect -67 -240 -63 -238
rect -35 -239 -32 -237
rect -14 -237 -8 -234
rect -14 -239 -11 -237
rect -86 -247 -77 -244
rect -113 -249 -104 -248
rect -108 -251 -104 -249
rect -86 -249 -83 -247
rect -95 -252 -83 -249
rect -95 -253 -92 -252
rect -105 -267 -102 -263
rect -86 -267 -83 -263
rect -54 -264 -51 -259
rect -23 -263 -20 -249
rect 1 -251 4 -194
rect 15 -204 18 -181
rect 53 -187 56 -180
rect 80 -178 83 -163
rect 71 -181 83 -178
rect 45 -190 56 -187
rect 53 -195 56 -190
rect 53 -198 57 -195
rect 15 -207 25 -204
rect 15 -228 18 -207
rect 53 -211 56 -206
rect 80 -204 83 -181
rect 87 -194 90 -153
rect 77 -207 83 -204
rect 45 -214 56 -211
rect 53 -219 56 -214
rect 53 -222 57 -219
rect 15 -231 25 -228
rect 53 -242 56 -230
rect 80 -228 83 -207
rect 87 -217 90 -198
rect 77 -231 83 -228
rect 87 -237 90 -221
rect 53 -245 59 -242
rect 1 -254 52 -251
rect -60 -267 -24 -264
rect -119 -270 -56 -267
rect 11 -273 14 -254
rect 39 -261 42 -254
rect 0 -276 14 -273
rect 49 -271 52 -254
rect 56 -253 59 -245
rect 56 -256 159 -253
rect 85 -264 151 -261
rect 85 -271 88 -264
rect 49 -274 88 -271
rect 11 -283 14 -276
rect 54 -281 57 -274
rect 72 -281 76 -274
rect 85 -287 88 -274
rect 120 -271 123 -264
rect 148 -283 151 -264
rect 156 -276 159 -256
rect 156 -279 219 -276
rect 148 -286 207 -283
rect 148 -293 151 -286
rect 179 -293 182 -286
rect 197 -293 201 -286
rect -268 -303 -205 -300
rect 2 -310 5 -303
rect 20 -310 23 -301
rect 64 -302 67 -301
rect 64 -305 76 -302
rect -268 -316 -257 -314
rect -5 -313 5 -310
rect 2 -315 5 -313
rect 13 -313 23 -310
rect 31 -311 55 -308
rect 20 -315 23 -313
rect 73 -314 76 -305
rect 94 -314 97 -307
rect -268 -317 -253 -316
rect -256 -324 -253 -317
rect -242 -319 -224 -315
rect 20 -318 32 -315
rect 41 -317 65 -314
rect 73 -317 86 -314
rect 29 -319 32 -318
rect 73 -319 76 -317
rect 94 -319 101 -314
rect -242 -324 -238 -319
rect -258 -327 -245 -324
rect -373 -351 -310 -348
rect -278 -351 -275 -344
rect -270 -345 -267 -342
rect -443 -359 -375 -356
rect -487 -362 -438 -359
rect -628 -372 -551 -368
rect -628 -445 -624 -372
rect -599 -381 -584 -378
rect -587 -388 -584 -381
rect -573 -388 -569 -372
rect -530 -374 -527 -367
rect -487 -369 -484 -362
rect -466 -369 -463 -362
rect -448 -369 -444 -362
rect -379 -364 -375 -359
rect -393 -366 -390 -364
rect -405 -369 -390 -366
rect -393 -372 -390 -369
rect -379 -367 -360 -364
rect -542 -377 -538 -374
rect -530 -377 -519 -374
rect -393 -376 -392 -372
rect -530 -379 -527 -377
rect -589 -391 -576 -388
rect -609 -415 -606 -408
rect -601 -409 -598 -406
rect -618 -417 -606 -415
rect -613 -418 -606 -417
rect -609 -421 -606 -418
rect -601 -421 -598 -414
rect -579 -415 -576 -391
rect -590 -419 -587 -416
rect -579 -418 -572 -415
rect -589 -432 -583 -428
rect -589 -434 -588 -432
rect -600 -437 -588 -434
rect -628 -449 -586 -445
rect -579 -446 -576 -418
rect -564 -424 -561 -408
rect -564 -426 -560 -424
rect -561 -429 -560 -426
rect -573 -435 -570 -430
rect -539 -435 -536 -389
rect -522 -394 -519 -377
rect -395 -377 -392 -376
rect -379 -376 -375 -367
rect -387 -377 -382 -376
rect -395 -379 -382 -377
rect -522 -397 -504 -394
rect -496 -396 -493 -387
rect -478 -396 -475 -389
rect -456 -390 -453 -389
rect -456 -393 -444 -390
rect -496 -399 -486 -396
rect -517 -403 -514 -400
rect -496 -401 -493 -399
rect -478 -399 -465 -396
rect -478 -401 -475 -399
rect -505 -404 -493 -401
rect -505 -405 -502 -404
rect -447 -402 -444 -393
rect -467 -406 -455 -403
rect -447 -403 -424 -402
rect -415 -403 -412 -396
rect -407 -397 -404 -394
rect -447 -405 -412 -403
rect -447 -407 -444 -405
rect -515 -419 -512 -415
rect -496 -419 -493 -415
rect -487 -418 -484 -411
rect -440 -415 -437 -405
rect -427 -406 -424 -405
rect -419 -406 -412 -405
rect -415 -409 -412 -406
rect -407 -409 -404 -402
rect -385 -403 -382 -379
rect -396 -407 -393 -404
rect -385 -406 -378 -403
rect -370 -412 -367 -396
rect -370 -414 -366 -412
rect -526 -422 -488 -419
rect -526 -435 -523 -422
rect -395 -420 -389 -416
rect -395 -422 -394 -420
rect -406 -425 -394 -422
rect -367 -417 -366 -414
rect -379 -423 -376 -418
rect -357 -423 -354 -351
rect -290 -353 -275 -351
rect -290 -354 -287 -353
rect -282 -354 -275 -353
rect -278 -357 -275 -354
rect -270 -357 -267 -350
rect -248 -351 -245 -327
rect -228 -324 -224 -319
rect -151 -323 -99 -320
rect -228 -325 -184 -324
rect -151 -325 -148 -323
rect -228 -328 -148 -325
rect -188 -341 -185 -328
rect -176 -335 -172 -328
rect -157 -335 -154 -328
rect -120 -330 -117 -323
rect -259 -355 -256 -352
rect -248 -354 -241 -351
rect -233 -360 -230 -344
rect -102 -354 -99 -323
rect 97 -323 101 -319
rect 118 -321 131 -318
rect 139 -320 142 -311
rect 157 -320 160 -313
rect 189 -314 192 -313
rect 189 -317 201 -314
rect 11 -333 14 -325
rect 20 -333 23 -329
rect 39 -333 42 -329
rect -11 -336 50 -333
rect -167 -356 -164 -355
rect -233 -362 -229 -360
rect -258 -368 -252 -364
rect -258 -370 -257 -368
rect -269 -373 -257 -370
rect -230 -365 -229 -362
rect -176 -359 -164 -356
rect -102 -357 -72 -354
rect -242 -371 -239 -366
rect -197 -368 -194 -361
rect -176 -368 -173 -359
rect -155 -365 -148 -362
rect -76 -366 -72 -357
rect -61 -356 -58 -354
rect -61 -359 -46 -356
rect -61 -366 -58 -359
rect -208 -371 -194 -368
rect -242 -374 -237 -371
rect -242 -378 -239 -374
rect -327 -381 -239 -378
rect -327 -413 -324 -381
rect -208 -393 -205 -371
rect -197 -373 -194 -371
rect -186 -371 -173 -368
rect -176 -373 -173 -371
rect -165 -372 -148 -369
rect -151 -379 -148 -372
rect -69 -369 -56 -366
rect -139 -379 -136 -370
rect -151 -382 -136 -379
rect -128 -380 -103 -377
rect -247 -396 -205 -393
rect -247 -410 -244 -396
rect -188 -398 -185 -383
rect -139 -384 -136 -382
rect -139 -387 -127 -384
rect -118 -387 -116 -383
rect -130 -388 -127 -387
rect -157 -398 -154 -393
rect -188 -401 -148 -398
rect -151 -402 -148 -401
rect -139 -402 -136 -398
rect -120 -402 -117 -398
rect -151 -405 -110 -402
rect -247 -413 -233 -410
rect -327 -416 -261 -413
rect -379 -426 -354 -423
rect -466 -431 -463 -427
rect -573 -438 -523 -435
rect -357 -432 -354 -426
rect -264 -428 -261 -416
rect -462 -435 -354 -432
rect -527 -441 -523 -438
rect -357 -441 -354 -435
rect -287 -431 -215 -428
rect -287 -441 -284 -431
rect -527 -444 -463 -441
rect -590 -522 -586 -449
rect -554 -449 -542 -446
rect -543 -451 -542 -449
rect -543 -455 -537 -451
rect -527 -453 -524 -444
rect -500 -448 -497 -444
rect -481 -448 -478 -444
rect -517 -453 -514 -451
rect -515 -457 -514 -453
rect -466 -449 -463 -444
rect -367 -444 -284 -441
rect -218 -438 -215 -431
rect -143 -438 -140 -405
rect -113 -413 -110 -405
rect -111 -418 -110 -413
rect -218 -441 -135 -438
rect -394 -449 -382 -446
rect -383 -451 -382 -449
rect -575 -466 -572 -465
rect -563 -465 -560 -462
rect -567 -466 -560 -465
rect -575 -468 -560 -466
rect -575 -508 -572 -468
rect -563 -475 -560 -468
rect -555 -469 -552 -462
rect -544 -467 -541 -464
rect -533 -468 -526 -465
rect -533 -472 -530 -468
rect -555 -477 -552 -474
rect -518 -475 -515 -457
rect -383 -455 -377 -451
rect -367 -453 -364 -444
rect -340 -448 -337 -444
rect -321 -448 -318 -444
rect -357 -453 -354 -451
rect -355 -457 -354 -453
rect -306 -449 -303 -444
rect -490 -459 -487 -458
rect -502 -463 -499 -460
rect -490 -460 -478 -459
rect -490 -462 -475 -460
rect -481 -463 -470 -462
rect -506 -469 -489 -466
rect -506 -472 -503 -469
rect -533 -492 -530 -477
rect -481 -476 -478 -463
rect -468 -473 -455 -470
rect -447 -471 -444 -469
rect -415 -466 -412 -465
rect -403 -465 -400 -462
rect -407 -466 -400 -465
rect -415 -468 -400 -466
rect -441 -471 -438 -468
rect -447 -474 -438 -471
rect -472 -480 -465 -477
rect -472 -484 -469 -480
rect -447 -483 -444 -474
rect -456 -486 -444 -483
rect -456 -487 -453 -486
rect -543 -495 -530 -492
rect -541 -502 -538 -495
rect -553 -505 -538 -502
rect -527 -504 -523 -495
rect -542 -509 -539 -505
rect -527 -507 -503 -504
rect -506 -522 -503 -507
rect -590 -523 -503 -522
rect -466 -514 -463 -507
rect -448 -514 -444 -507
rect -415 -508 -412 -468
rect -403 -475 -400 -468
rect -395 -469 -392 -462
rect -384 -467 -381 -464
rect -373 -468 -366 -465
rect -373 -472 -370 -468
rect -395 -477 -392 -474
rect -358 -475 -355 -457
rect -330 -459 -327 -458
rect -342 -463 -339 -460
rect -330 -460 -318 -459
rect -330 -462 -315 -460
rect -321 -463 -310 -462
rect -346 -469 -329 -466
rect -346 -472 -343 -469
rect -373 -492 -370 -477
rect -321 -476 -318 -463
rect -308 -473 -295 -470
rect -287 -471 -284 -469
rect -281 -471 -278 -441
rect -245 -446 -233 -443
rect -234 -448 -233 -446
rect -234 -452 -228 -448
rect -218 -450 -215 -441
rect -191 -445 -188 -441
rect -172 -445 -169 -441
rect -208 -450 -205 -448
rect -206 -454 -205 -450
rect -157 -446 -154 -441
rect -287 -474 -278 -471
rect -266 -463 -263 -462
rect -254 -462 -251 -459
rect -258 -463 -251 -462
rect -266 -465 -251 -463
rect -312 -480 -305 -477
rect -312 -484 -309 -480
rect -287 -483 -284 -474
rect -296 -486 -284 -483
rect -296 -487 -293 -486
rect -383 -495 -370 -492
rect -381 -502 -378 -495
rect -393 -505 -378 -502
rect -367 -504 -363 -495
rect -382 -508 -379 -505
rect -367 -507 -343 -504
rect -500 -523 -497 -516
rect -476 -517 -438 -514
rect -476 -522 -472 -517
rect -346 -522 -343 -507
rect -266 -504 -263 -465
rect -254 -472 -251 -465
rect -246 -466 -243 -459
rect -235 -464 -232 -461
rect -224 -465 -217 -462
rect -224 -469 -221 -465
rect -246 -474 -243 -471
rect -209 -472 -206 -454
rect -181 -456 -178 -455
rect -193 -460 -190 -457
rect -181 -457 -169 -456
rect -181 -459 -166 -457
rect -172 -460 -161 -459
rect -197 -466 -180 -463
rect -197 -469 -194 -466
rect -224 -489 -221 -474
rect -172 -473 -169 -460
rect -159 -470 -146 -467
rect -138 -468 -135 -466
rect -132 -467 -129 -431
rect -113 -435 -110 -418
rect -106 -429 -103 -380
rect -84 -402 -81 -386
rect -69 -391 -66 -369
rect -47 -387 -44 -384
rect -73 -396 -72 -393
rect -67 -396 -66 -391
rect -58 -397 -55 -394
rect -47 -399 -44 -392
rect -85 -404 -81 -402
rect -39 -393 -36 -386
rect -27 -393 -24 -360
rect -39 -395 -24 -393
rect -11 -394 -8 -336
rect 47 -344 50 -336
rect 54 -344 57 -339
rect 85 -343 88 -329
rect 98 -332 101 -323
rect 139 -323 149 -320
rect 113 -326 121 -325
rect 118 -328 121 -326
rect 139 -325 142 -323
rect 157 -323 180 -320
rect 157 -325 160 -323
rect 130 -328 142 -325
rect 130 -329 133 -328
rect 198 -326 201 -317
rect 99 -337 101 -332
rect 166 -330 190 -327
rect 198 -329 211 -326
rect 166 -331 170 -330
rect 198 -331 201 -329
rect 120 -343 123 -339
rect 139 -343 142 -339
rect 148 -343 151 -335
rect 85 -344 176 -343
rect 47 -346 176 -344
rect 47 -347 88 -346
rect -39 -396 -32 -395
rect -39 -399 -36 -396
rect -27 -396 -24 -395
rect -21 -397 -8 -394
rect 91 -363 94 -361
rect 91 -366 101 -363
rect 91 -396 94 -366
rect 148 -374 151 -349
rect 173 -356 176 -346
rect 208 -349 211 -329
rect 179 -356 182 -351
rect 173 -359 204 -356
rect 154 -364 157 -359
rect 173 -363 176 -359
rect 216 -363 219 -279
rect 169 -366 176 -363
rect 155 -376 159 -373
rect 155 -382 158 -376
rect 141 -385 158 -382
rect 173 -382 176 -366
rect 169 -385 176 -382
rect 181 -366 219 -363
rect 150 -393 153 -385
rect 181 -389 184 -366
rect 133 -396 153 -393
rect 158 -392 184 -389
rect -85 -407 -84 -404
rect -75 -413 -72 -408
rect -94 -416 -72 -413
rect -62 -410 -56 -406
rect -57 -412 -56 -410
rect -57 -415 -45 -412
rect -21 -422 -18 -397
rect 43 -399 111 -396
rect 49 -406 52 -399
rect 67 -406 71 -399
rect 83 -406 86 -399
rect 101 -406 105 -399
rect 158 -400 161 -392
rect 118 -403 161 -400
rect -21 -425 -2 -422
rect -106 -432 -14 -429
rect -113 -438 -63 -435
rect -5 -438 -2 -425
rect 59 -427 62 -426
rect 93 -427 96 -426
rect 59 -430 71 -427
rect 93 -430 105 -427
rect -66 -441 4 -438
rect -93 -446 -81 -443
rect -82 -448 -81 -446
rect -82 -452 -76 -448
rect -66 -450 -63 -441
rect -39 -445 -36 -441
rect -20 -445 -17 -441
rect -56 -450 -53 -448
rect -54 -454 -53 -450
rect -5 -446 -2 -441
rect -114 -463 -111 -462
rect -102 -462 -99 -459
rect -106 -463 -99 -462
rect -114 -465 -99 -463
rect -138 -471 -132 -468
rect -163 -477 -156 -474
rect -163 -481 -160 -477
rect -138 -480 -135 -471
rect -147 -483 -135 -480
rect -147 -484 -144 -483
rect -234 -492 -221 -489
rect -232 -499 -229 -492
rect -244 -502 -229 -499
rect -218 -501 -214 -492
rect -476 -523 -343 -522
rect -306 -514 -303 -507
rect -288 -514 -284 -507
rect -233 -506 -230 -502
rect -218 -504 -194 -501
rect -197 -514 -194 -504
rect -114 -503 -111 -465
rect -102 -472 -99 -465
rect -94 -466 -91 -459
rect -83 -464 -80 -461
rect -72 -465 -65 -462
rect -72 -469 -69 -465
rect -94 -474 -91 -471
rect -57 -472 -54 -454
rect -29 -456 -26 -455
rect -41 -460 -38 -457
rect -29 -457 -17 -456
rect -29 -459 -14 -457
rect -20 -460 -9 -459
rect -45 -466 -28 -463
rect -45 -469 -42 -466
rect -72 -489 -69 -474
rect -20 -473 -17 -460
rect -7 -470 6 -467
rect 14 -468 17 -466
rect 20 -468 23 -434
rect 44 -436 50 -433
rect 14 -471 23 -468
rect 36 -443 60 -440
rect 68 -440 71 -430
rect 82 -437 84 -433
rect 102 -439 105 -430
rect 118 -439 121 -403
rect 68 -443 94 -440
rect 102 -442 121 -439
rect -11 -477 -4 -474
rect -11 -481 -8 -477
rect 14 -480 17 -471
rect 5 -483 17 -480
rect 5 -484 8 -483
rect -82 -492 -69 -489
rect -80 -499 -77 -492
rect -92 -502 -77 -499
rect -82 -503 -77 -502
rect -340 -523 -337 -516
rect -316 -517 -194 -514
rect -316 -523 -312 -517
rect -197 -520 -194 -517
rect -157 -511 -154 -504
rect -139 -511 -135 -504
rect -66 -501 -62 -492
rect 36 -495 39 -443
rect 68 -444 71 -443
rect 102 -444 105 -442
rect 49 -468 52 -464
rect 47 -469 52 -468
rect 83 -469 86 -464
rect 47 -472 108 -469
rect -66 -504 -42 -501
rect -45 -511 -42 -504
rect -191 -520 -188 -513
rect -167 -514 -42 -511
rect -167 -520 -163 -514
rect -197 -523 -163 -520
rect -45 -520 -42 -514
rect -5 -511 -2 -504
rect 13 -511 17 -504
rect -39 -520 -36 -513
rect -15 -514 23 -511
rect -15 -520 -11 -514
rect -45 -523 -11 -520
rect -590 -526 -312 -523
rect -618 -553 -615 -541
rect -580 -544 -575 -543
rect -588 -548 -572 -544
rect -618 -556 -608 -553
rect -618 -578 -615 -556
rect -580 -560 -577 -555
rect -562 -556 -550 -553
rect -591 -563 -576 -560
rect -591 -569 -588 -563
rect -618 -581 -608 -578
rect -618 -603 -615 -581
rect -580 -585 -577 -580
rect -553 -578 -550 -556
rect -539 -554 -536 -542
rect -509 -549 -493 -545
rect -457 -551 -454 -539
rect -427 -546 -411 -542
rect -539 -557 -529 -554
rect -556 -581 -550 -578
rect -591 -588 -576 -585
rect -591 -594 -588 -588
rect -618 -606 -608 -603
rect -618 -621 -615 -606
rect -580 -612 -577 -605
rect -553 -603 -550 -581
rect -546 -592 -543 -571
rect -556 -606 -550 -603
rect -588 -616 -572 -612
rect -618 -624 -608 -621
rect -618 -647 -615 -624
rect -580 -630 -577 -623
rect -553 -621 -550 -606
rect -562 -624 -550 -621
rect -588 -633 -577 -630
rect -580 -638 -577 -633
rect -580 -641 -576 -638
rect -618 -650 -608 -647
rect -618 -671 -615 -650
rect -580 -654 -577 -649
rect -553 -647 -550 -624
rect -546 -637 -543 -596
rect -556 -650 -550 -647
rect -588 -657 -577 -654
rect -580 -662 -577 -657
rect -580 -665 -576 -662
rect -618 -674 -608 -671
rect -618 -680 -615 -674
rect -580 -680 -577 -673
rect -553 -671 -550 -650
rect -546 -660 -543 -641
rect -556 -674 -550 -671
rect -547 -673 -543 -664
rect -539 -579 -536 -557
rect -501 -561 -498 -556
rect -457 -554 -447 -551
rect -483 -557 -471 -554
rect -512 -564 -497 -561
rect -512 -570 -509 -564
rect -539 -582 -529 -579
rect -539 -604 -536 -582
rect -501 -586 -498 -581
rect -474 -579 -471 -557
rect -477 -582 -471 -579
rect -512 -589 -497 -586
rect -512 -595 -509 -589
rect -539 -607 -529 -604
rect -539 -622 -536 -607
rect -501 -613 -498 -606
rect -474 -604 -471 -582
rect -467 -593 -464 -572
rect -477 -607 -471 -604
rect -509 -617 -493 -613
rect -539 -625 -529 -622
rect -539 -648 -536 -625
rect -501 -631 -498 -624
rect -474 -622 -471 -607
rect -483 -625 -471 -622
rect -509 -634 -498 -631
rect -501 -639 -498 -634
rect -501 -642 -497 -639
rect -539 -651 -529 -648
rect -539 -672 -536 -651
rect -501 -655 -498 -650
rect -474 -648 -471 -625
rect -467 -638 -464 -597
rect -477 -651 -471 -648
rect -509 -658 -498 -655
rect -501 -663 -498 -658
rect -501 -666 -497 -663
rect -539 -675 -529 -672
rect -501 -681 -498 -674
rect -474 -672 -471 -651
rect -467 -661 -464 -642
rect -477 -675 -471 -672
rect -467 -675 -464 -665
rect -457 -576 -454 -554
rect -419 -558 -416 -553
rect -401 -554 -389 -551
rect -430 -561 -415 -558
rect -430 -567 -427 -561
rect -457 -579 -447 -576
rect -457 -601 -454 -579
rect -419 -583 -416 -578
rect -392 -576 -389 -554
rect -373 -552 -370 -540
rect -343 -547 -327 -543
rect -373 -555 -363 -552
rect -291 -551 -288 -539
rect -261 -546 -245 -542
rect -395 -579 -389 -576
rect -430 -586 -415 -583
rect -430 -592 -427 -586
rect -457 -604 -447 -601
rect -457 -619 -454 -604
rect -419 -610 -416 -603
rect -392 -601 -389 -579
rect -385 -590 -382 -569
rect -395 -604 -389 -601
rect -427 -614 -411 -610
rect -457 -622 -447 -619
rect -457 -645 -454 -622
rect -419 -628 -416 -621
rect -392 -619 -389 -604
rect -401 -622 -389 -619
rect -427 -631 -416 -628
rect -419 -636 -416 -631
rect -419 -639 -415 -636
rect -457 -648 -447 -645
rect -457 -669 -454 -648
rect -419 -652 -416 -647
rect -392 -645 -389 -622
rect -385 -635 -382 -594
rect -395 -648 -389 -645
rect -427 -655 -416 -652
rect -419 -660 -416 -655
rect -419 -663 -415 -660
rect -457 -672 -447 -669
rect -457 -686 -454 -672
rect -419 -678 -416 -671
rect -392 -669 -389 -648
rect -385 -658 -382 -639
rect -395 -672 -389 -669
rect -385 -674 -382 -662
rect -373 -577 -370 -555
rect -335 -559 -332 -554
rect -317 -555 -305 -552
rect -346 -562 -331 -559
rect -346 -568 -343 -562
rect -373 -580 -363 -577
rect -373 -602 -370 -580
rect -335 -584 -332 -579
rect -308 -577 -305 -555
rect -291 -554 -281 -551
rect -311 -580 -305 -577
rect -346 -587 -331 -584
rect -346 -593 -343 -587
rect -373 -605 -363 -602
rect -373 -620 -370 -605
rect -335 -611 -332 -604
rect -308 -602 -305 -580
rect -301 -591 -298 -570
rect -311 -605 -305 -602
rect -343 -615 -327 -611
rect -373 -623 -363 -620
rect -373 -646 -370 -623
rect -335 -629 -332 -622
rect -308 -620 -305 -605
rect -317 -623 -305 -620
rect -343 -632 -332 -629
rect -335 -637 -332 -632
rect -335 -640 -331 -637
rect -373 -649 -363 -646
rect -373 -670 -370 -649
rect -335 -653 -332 -648
rect -308 -646 -305 -623
rect -301 -636 -298 -595
rect -311 -649 -305 -646
rect -343 -656 -332 -653
rect -335 -661 -332 -656
rect -335 -664 -331 -661
rect -373 -673 -363 -670
rect -373 -682 -370 -673
rect -335 -679 -332 -672
rect -308 -670 -305 -649
rect -301 -659 -298 -640
rect -311 -673 -305 -670
rect -301 -675 -298 -663
rect -291 -576 -288 -554
rect -253 -558 -250 -553
rect -205 -551 -202 -539
rect -175 -546 -159 -542
rect -235 -554 -223 -551
rect -264 -561 -249 -558
rect -264 -567 -261 -561
rect -291 -579 -281 -576
rect -291 -601 -288 -579
rect -253 -583 -250 -578
rect -226 -576 -223 -554
rect -205 -554 -195 -551
rect -229 -579 -223 -576
rect -264 -586 -249 -583
rect -264 -592 -261 -586
rect -291 -604 -281 -601
rect -291 -619 -288 -604
rect -253 -610 -250 -603
rect -226 -601 -223 -579
rect -219 -590 -216 -569
rect -229 -604 -223 -601
rect -261 -614 -245 -610
rect -291 -622 -281 -619
rect -291 -645 -288 -622
rect -253 -628 -250 -621
rect -226 -619 -223 -604
rect -235 -622 -223 -619
rect -261 -631 -250 -628
rect -253 -636 -250 -631
rect -253 -639 -249 -636
rect -291 -648 -281 -645
rect -291 -669 -288 -648
rect -253 -652 -250 -647
rect -226 -645 -223 -622
rect -219 -635 -216 -594
rect -229 -648 -223 -645
rect -261 -655 -250 -652
rect -253 -660 -250 -655
rect -253 -663 -249 -660
rect -291 -672 -281 -669
rect -291 -682 -288 -672
rect -253 -678 -250 -671
rect -226 -669 -223 -648
rect -219 -658 -216 -639
rect -229 -672 -223 -669
rect -219 -675 -216 -662
rect -205 -576 -202 -554
rect -167 -558 -164 -553
rect -149 -554 -137 -551
rect -178 -561 -163 -558
rect -178 -567 -175 -561
rect -205 -579 -195 -576
rect -205 -601 -202 -579
rect -167 -583 -164 -578
rect -140 -576 -137 -554
rect -120 -552 -117 -540
rect -90 -547 -74 -543
rect -120 -555 -110 -552
rect -143 -579 -137 -576
rect -178 -586 -163 -583
rect -178 -592 -175 -586
rect -205 -604 -195 -601
rect -205 -619 -202 -604
rect -167 -610 -164 -603
rect -140 -601 -137 -579
rect -133 -590 -130 -569
rect -143 -604 -137 -601
rect -175 -614 -159 -610
rect -205 -622 -195 -619
rect -205 -645 -202 -622
rect -167 -628 -164 -621
rect -140 -619 -137 -604
rect -149 -622 -137 -619
rect -175 -631 -164 -628
rect -167 -636 -164 -631
rect -167 -639 -163 -636
rect -205 -648 -195 -645
rect -205 -669 -202 -648
rect -167 -652 -164 -647
rect -140 -645 -137 -622
rect -133 -635 -130 -594
rect -143 -648 -137 -645
rect -175 -655 -164 -652
rect -167 -660 -164 -655
rect -167 -663 -163 -660
rect -205 -672 -195 -669
rect -205 -682 -202 -672
rect -167 -678 -164 -671
rect -140 -669 -137 -648
rect -133 -658 -130 -639
rect -143 -672 -137 -669
rect -133 -675 -130 -662
rect -120 -577 -117 -555
rect -82 -559 -79 -554
rect -37 -552 -34 -540
rect -7 -544 0 -543
rect 5 -544 9 -543
rect -7 -547 9 -544
rect -64 -555 -52 -552
rect -93 -562 -78 -559
rect -93 -568 -90 -562
rect -120 -580 -110 -577
rect -120 -602 -117 -580
rect -82 -584 -79 -579
rect -55 -577 -52 -555
rect -37 -555 -27 -552
rect -58 -580 -52 -577
rect -93 -587 -78 -584
rect -93 -593 -90 -587
rect -120 -605 -110 -602
rect -120 -620 -117 -605
rect -82 -611 -79 -604
rect -55 -602 -52 -580
rect -48 -591 -45 -570
rect -58 -605 -52 -602
rect -90 -615 -74 -611
rect -120 -623 -110 -620
rect -120 -646 -117 -623
rect -82 -629 -79 -622
rect -55 -620 -52 -605
rect -64 -623 -52 -620
rect -90 -632 -79 -629
rect -82 -637 -79 -632
rect -82 -640 -78 -637
rect -120 -649 -110 -646
rect -120 -670 -117 -649
rect -82 -653 -79 -648
rect -55 -646 -52 -623
rect -48 -636 -45 -595
rect -58 -649 -52 -646
rect -90 -656 -79 -653
rect -82 -661 -79 -656
rect -82 -664 -78 -661
rect -120 -673 -110 -670
rect -82 -679 -79 -672
rect -55 -670 -52 -649
rect -48 -659 -45 -640
rect -58 -673 -52 -670
rect -48 -675 -45 -663
rect -37 -577 -34 -555
rect 1 -559 4 -554
rect 47 -552 50 -540
rect 77 -547 93 -543
rect 19 -555 31 -552
rect -10 -562 5 -559
rect -10 -568 -7 -562
rect -37 -580 -27 -577
rect -37 -602 -34 -580
rect 1 -584 4 -579
rect 28 -577 31 -555
rect 47 -555 57 -552
rect 25 -580 31 -577
rect -10 -587 5 -584
rect -10 -593 -7 -587
rect -37 -605 -27 -602
rect -37 -620 -34 -605
rect 1 -611 4 -604
rect 28 -602 31 -580
rect 35 -591 38 -570
rect 25 -605 31 -602
rect -7 -615 9 -611
rect -37 -623 -27 -620
rect -37 -646 -34 -623
rect 1 -629 4 -622
rect 28 -620 31 -605
rect 19 -623 31 -620
rect -7 -632 4 -629
rect 1 -637 4 -632
rect 1 -640 5 -637
rect -37 -649 -27 -646
rect -37 -670 -34 -649
rect 1 -653 4 -648
rect 28 -646 31 -623
rect 35 -636 38 -595
rect 25 -649 31 -646
rect -7 -656 4 -653
rect 1 -661 4 -656
rect 1 -664 5 -661
rect -37 -673 -27 -670
rect -37 -682 -34 -673
rect 1 -679 4 -672
rect 28 -670 31 -649
rect 35 -659 38 -640
rect 25 -673 31 -670
rect 35 -675 38 -663
rect 47 -577 50 -555
rect 85 -559 88 -554
rect 103 -555 115 -552
rect 74 -562 89 -559
rect 74 -568 77 -562
rect 47 -580 57 -577
rect 47 -602 50 -580
rect 85 -584 88 -579
rect 112 -577 115 -555
rect 109 -580 115 -577
rect 74 -587 89 -584
rect 74 -593 77 -587
rect 47 -605 57 -602
rect 47 -620 50 -605
rect 85 -611 88 -604
rect 112 -602 115 -580
rect 119 -591 122 -570
rect 109 -605 115 -602
rect 77 -615 93 -611
rect 47 -623 57 -620
rect 47 -646 50 -623
rect 85 -629 88 -622
rect 112 -620 115 -605
rect 103 -623 115 -620
rect 77 -632 88 -629
rect 85 -637 88 -632
rect 85 -640 89 -637
rect 47 -649 57 -646
rect 47 -670 50 -649
rect 85 -653 88 -648
rect 112 -646 115 -623
rect 119 -636 122 -595
rect 109 -649 115 -646
rect 77 -656 88 -653
rect 85 -661 88 -656
rect 85 -664 89 -661
rect 47 -673 57 -670
rect 47 -682 50 -673
rect 85 -679 88 -672
rect 112 -670 115 -649
rect 119 -659 122 -640
rect 109 -673 115 -670
rect 119 -675 122 -663
<< m2contact >>
rect -91 -108 -85 -103
rect -124 -140 -119 -135
rect -294 -196 -289 -191
rect -310 -221 -305 -216
rect -105 -149 -100 -144
rect -121 -192 -116 -187
rect -50 -186 -45 -181
rect -329 -230 -324 -225
rect -384 -267 -379 -262
rect -496 -316 -491 -311
rect -596 -355 -591 -349
rect -218 -281 -213 -276
rect -426 -320 -421 -315
rect -322 -326 -317 -321
rect -8 -239 -3 -234
rect -257 -316 -252 -311
rect -271 -350 -266 -345
rect -602 -414 -597 -409
rect -588 -437 -583 -432
rect -560 -429 -555 -424
rect -392 -377 -387 -372
rect -408 -402 -403 -397
rect -488 -423 -483 -418
rect -394 -425 -389 -420
rect -366 -417 -361 -412
rect -257 -373 -252 -368
rect -229 -365 -224 -360
rect -233 -413 -228 -408
rect -467 -436 -462 -431
rect -580 -451 -575 -446
rect -542 -451 -537 -446
rect -514 -454 -509 -449
rect -281 -441 -276 -435
rect -116 -418 -111 -413
rect -133 -431 -128 -426
rect -382 -451 -377 -446
rect -556 -474 -551 -469
rect -534 -477 -529 -472
rect -354 -454 -349 -449
rect -475 -462 -470 -457
rect -507 -477 -502 -472
rect -473 -474 -468 -469
rect -576 -513 -571 -508
rect -543 -514 -538 -509
rect -396 -474 -391 -469
rect -374 -477 -369 -472
rect -315 -462 -310 -457
rect -347 -477 -342 -472
rect -313 -474 -308 -469
rect -233 -448 -228 -443
rect -205 -451 -200 -446
rect -416 -513 -411 -508
rect -383 -513 -378 -508
rect -247 -471 -242 -466
rect -225 -474 -220 -469
rect -198 -474 -193 -469
rect -164 -471 -159 -466
rect -72 -396 -67 -391
rect -48 -392 -43 -387
rect -90 -407 -85 -402
rect 113 -331 118 -326
rect 94 -337 99 -332
rect 143 -354 148 -349
rect 154 -359 159 -354
rect 208 -354 213 -349
rect 128 -396 133 -391
rect -99 -417 -94 -412
rect -62 -415 -57 -410
rect -14 -433 -9 -428
rect -81 -448 -76 -443
rect -53 -451 -48 -446
rect 4 -442 9 -437
rect -267 -509 -262 -504
rect -234 -511 -229 -506
rect -95 -471 -90 -466
rect -73 -474 -68 -469
rect -14 -459 -9 -454
rect -46 -474 -41 -469
rect -12 -471 -7 -466
rect 39 -437 44 -432
rect 77 -437 82 -432
rect -115 -508 -110 -503
rect -82 -508 -77 -503
rect 42 -473 47 -468
rect 36 -500 41 -495
rect -580 -543 -575 -538
rect -502 -545 -497 -540
rect -420 -542 -415 -537
rect -547 -678 -542 -673
rect -336 -543 -331 -538
rect -254 -542 -249 -537
rect -468 -681 -462 -675
rect -386 -679 -381 -674
rect -168 -542 -163 -537
rect -302 -680 -297 -675
rect -220 -680 -215 -675
rect 0 -544 5 -539
rect -134 -680 -129 -675
rect 84 -543 89 -538
rect -49 -680 -44 -675
rect 34 -680 39 -675
rect 118 -680 123 -675
<< metal2 >>
rect -90 -121 -87 -108
rect -119 -139 -102 -136
rect -105 -144 -102 -139
rect -112 -185 -50 -182
rect -293 -201 -290 -196
rect -327 -220 -310 -217
rect -327 -225 -324 -220
rect -119 -223 -116 -192
rect -238 -228 -227 -225
rect -434 -234 -431 -233
rect -496 -237 -431 -234
rect -496 -311 -493 -237
rect -621 -355 -596 -352
rect -621 -410 -618 -355
rect -434 -398 -431 -237
rect -238 -245 -235 -228
rect -203 -226 -116 -223
rect -320 -248 -235 -245
rect -320 -263 -317 -248
rect -379 -266 -317 -263
rect -425 -281 -366 -278
rect -425 -315 -422 -281
rect -320 -321 -317 -266
rect -311 -316 -308 -267
rect -217 -308 -214 -281
rect -256 -311 -214 -308
rect -311 -319 -298 -316
rect -317 -326 -306 -323
rect -309 -352 -306 -326
rect -352 -355 -306 -352
rect -393 -377 -392 -374
rect -387 -377 -383 -374
rect -386 -381 -383 -377
rect -434 -401 -408 -398
rect -621 -413 -602 -410
rect -617 -449 -614 -422
rect -586 -439 -583 -437
rect -559 -439 -556 -429
rect -586 -442 -556 -439
rect -522 -439 -519 -405
rect -483 -422 -467 -419
rect -470 -435 -467 -422
rect -392 -427 -389 -425
rect -365 -427 -362 -417
rect -392 -430 -362 -427
rect -352 -436 -349 -355
rect -301 -359 -298 -319
rect -293 -346 -289 -313
rect -203 -317 -200 -226
rect -112 -240 -109 -185
rect -63 -200 -4 -197
rect -7 -234 -4 -200
rect -220 -320 -200 -317
rect -2 -289 102 -286
rect -293 -349 -271 -346
rect -345 -362 -298 -359
rect -345 -428 -342 -362
rect -286 -368 -283 -358
rect -335 -371 -283 -368
rect -335 -420 -332 -371
rect -255 -375 -252 -373
rect -228 -375 -225 -365
rect -255 -378 -225 -375
rect -220 -383 -217 -320
rect -321 -386 -217 -383
rect -321 -408 -318 -386
rect -99 -396 -72 -393
rect -17 -388 -14 -346
rect -43 -391 -14 -388
rect -99 -403 -96 -396
rect -124 -406 -96 -403
rect -321 -411 -256 -408
rect -335 -423 -267 -420
rect -345 -431 -277 -428
rect -280 -435 -277 -431
rect -352 -439 -311 -436
rect -522 -442 -471 -439
rect -617 -452 -591 -449
rect -537 -451 -514 -450
rect -594 -496 -591 -452
rect -579 -470 -576 -451
rect -541 -453 -514 -451
rect -474 -457 -471 -442
rect -579 -473 -556 -470
rect -506 -470 -503 -468
rect -506 -472 -473 -470
rect -529 -476 -507 -473
rect -502 -473 -473 -472
rect -419 -470 -416 -450
rect -377 -451 -354 -450
rect -381 -453 -354 -451
rect -314 -457 -311 -439
rect -270 -467 -267 -423
rect -259 -423 -256 -411
rect -228 -412 -197 -409
rect -259 -426 -208 -423
rect -124 -424 -121 -406
rect -2 -403 1 -289
rect 99 -325 102 -289
rect 99 -328 106 -325
rect 103 -337 106 -328
rect 113 -337 116 -331
rect 95 -348 98 -337
rect 103 -340 116 -337
rect 95 -349 148 -348
rect 95 -351 143 -349
rect 154 -353 208 -350
rect 154 -354 159 -353
rect 31 -397 42 -394
rect -13 -406 1 -403
rect -111 -416 -99 -413
rect -89 -417 -86 -407
rect -62 -417 -59 -415
rect -89 -420 -59 -417
rect -211 -427 -208 -426
rect -211 -430 -133 -427
rect -124 -427 -115 -424
rect -228 -448 -205 -447
rect -232 -450 -205 -448
rect -419 -473 -396 -470
rect -346 -470 -343 -468
rect -346 -472 -313 -470
rect -369 -476 -347 -473
rect -342 -473 -313 -472
rect -270 -470 -247 -467
rect -197 -467 -194 -465
rect -197 -469 -164 -467
rect -220 -473 -198 -470
rect -193 -470 -164 -469
rect -118 -467 -115 -427
rect -13 -428 -10 -406
rect -76 -448 -53 -447
rect -80 -450 -53 -448
rect -13 -454 -10 -433
rect 39 -432 42 -397
rect 78 -395 128 -392
rect 78 -432 81 -395
rect 9 -441 27 -438
rect -118 -470 -95 -467
rect -45 -467 -42 -465
rect -45 -469 -12 -467
rect -68 -473 -46 -470
rect -41 -470 -12 -469
rect 24 -469 27 -441
rect 24 -472 42 -469
rect -628 -499 36 -496
rect -628 -536 -625 -499
rect -575 -529 -572 -513
rect -575 -532 -552 -529
rect -628 -538 -577 -536
rect -628 -539 -580 -538
rect -555 -540 -552 -532
rect -542 -532 -539 -514
rect -415 -525 -412 -513
rect -382 -525 -379 -513
rect -266 -517 -263 -509
rect -266 -520 -239 -517
rect -415 -528 -388 -525
rect -382 -528 -250 -525
rect -391 -532 -388 -528
rect -542 -535 -454 -532
rect -391 -535 -332 -532
rect -457 -538 -454 -535
rect -555 -543 -502 -540
rect -457 -541 -420 -538
rect -336 -538 -332 -535
rect -253 -537 -250 -528
rect -242 -528 -239 -520
rect -233 -521 -230 -511
rect -233 -524 -138 -521
rect -242 -531 -165 -528
rect -168 -537 -165 -531
rect -114 -531 -110 -508
rect -81 -523 -78 -508
rect -81 -526 88 -523
rect -114 -534 4 -531
rect 0 -539 4 -534
rect 85 -538 88 -526
rect -542 -678 -468 -675
rect -462 -678 -386 -675
rect -381 -678 -302 -675
rect -297 -678 -220 -675
rect -215 -678 -134 -675
rect -129 -678 -49 -675
rect -44 -678 34 -675
rect 39 -678 118 -675
<< m3contact >>
rect -366 -282 -361 -277
rect -68 -201 -63 -196
rect -197 -413 -192 -408
rect 26 -398 31 -393
rect -138 -525 -133 -520
rect -458 -687 -453 -682
<< m123contact >>
rect -23 -176 -18 -171
rect -41 -181 -36 -176
rect -215 -201 -210 -196
rect -165 -205 -160 -200
rect -443 -265 -438 -260
rect -547 -378 -542 -373
rect -411 -257 -406 -252
rect -372 -321 -367 -316
rect -312 -267 -307 -262
rect -269 -286 -264 -281
rect -321 -337 -316 -332
rect -410 -349 -405 -344
rect -522 -405 -517 -400
rect -618 -422 -613 -417
rect -587 -420 -582 -415
rect -472 -408 -467 -403
rect -424 -410 -419 -405
rect -393 -408 -388 -403
rect -441 -420 -436 -415
rect -112 -245 -107 -240
rect -68 -245 -63 -240
rect -113 -254 -108 -249
rect -24 -268 -19 -263
rect -5 -276 0 -271
rect -287 -358 -282 -353
rect -256 -356 -251 -351
rect -27 -360 -22 -355
rect -116 -388 -111 -383
rect -63 -398 -58 -393
rect -32 -400 -27 -395
rect -572 -466 -567 -461
rect -507 -463 -502 -458
rect -541 -468 -536 -463
rect -441 -468 -436 -463
rect -412 -466 -407 -461
rect -347 -463 -342 -458
rect -381 -468 -376 -463
rect 113 -322 118 -317
rect 165 -336 170 -331
rect 89 -361 94 -356
rect -263 -463 -258 -458
rect -198 -460 -193 -455
rect -166 -459 -161 -454
rect -232 -465 -227 -460
rect 19 -434 24 -429
rect -111 -463 -106 -458
rect -46 -460 -41 -455
rect -80 -465 -75 -460
rect -132 -472 -127 -467
rect -473 -489 -468 -484
rect -313 -489 -308 -484
rect -164 -486 -159 -481
rect -12 -486 -7 -481
rect -83 -543 -78 -538
rect -619 -685 -614 -680
rect -540 -687 -535 -682
rect -374 -687 -369 -682
rect -292 -687 -287 -682
rect -206 -687 -201 -682
rect -121 -687 -116 -682
rect -38 -687 -33 -682
rect 46 -687 51 -682
<< metal3 >>
rect -230 -181 -41 -178
rect -230 -210 -227 -181
rect -69 -196 -62 -195
rect -69 -197 -68 -196
rect -161 -200 -68 -197
rect -311 -213 -227 -210
rect -214 -212 -211 -201
rect -160 -203 -158 -200
rect -69 -201 -68 -200
rect -63 -201 -62 -196
rect -69 -202 -62 -201
rect -546 -325 -491 -322
rect -546 -373 -543 -325
rect -494 -326 -491 -325
rect -494 -329 -470 -326
rect -522 -334 -506 -331
rect -586 -377 -547 -374
rect -586 -415 -583 -377
rect -522 -400 -519 -334
rect -441 -353 -438 -265
rect -410 -344 -407 -257
rect -311 -262 -308 -213
rect -197 -232 -122 -229
rect -367 -277 -360 -276
rect -367 -282 -366 -277
rect -361 -278 -360 -277
rect -361 -281 -268 -278
rect -361 -282 -360 -281
rect -367 -283 -360 -282
rect -271 -284 -269 -281
rect -367 -321 -365 -316
rect -368 -334 -365 -321
rect -197 -324 -194 -232
rect -184 -315 -181 -232
rect -125 -241 -122 -232
rect -125 -244 -112 -241
rect -129 -252 -113 -249
rect -67 -271 -64 -245
rect -22 -263 -19 -176
rect -131 -274 -64 -271
rect -184 -318 -104 -315
rect -214 -327 -194 -324
rect -368 -337 -357 -334
rect -365 -338 -362 -337
rect -471 -356 -438 -353
rect -471 -403 -468 -356
rect -321 -354 -317 -337
rect -285 -353 -256 -352
rect -393 -358 -317 -354
rect -282 -355 -256 -353
rect -214 -389 -211 -327
rect -107 -384 -104 -318
rect -4 -329 -1 -276
rect 107 -322 113 -318
rect -4 -332 10 -329
rect 7 -338 10 -332
rect 7 -341 46 -338
rect -31 -351 -24 -348
rect -27 -355 -24 -351
rect -6 -349 35 -346
rect -111 -387 -104 -384
rect -313 -392 -211 -389
rect -313 -402 -310 -392
rect -58 -395 -29 -394
rect -58 -397 -32 -395
rect -6 -398 -3 -349
rect -17 -401 -3 -398
rect 2 -354 10 -353
rect -422 -405 -393 -404
rect -616 -417 -587 -416
rect -613 -419 -587 -417
rect -544 -463 -507 -460
rect -471 -463 -468 -408
rect -419 -407 -393 -405
rect -313 -405 -249 -402
rect -252 -415 -249 -405
rect -192 -412 -186 -409
rect -436 -420 -432 -416
rect -252 -418 -201 -415
rect -435 -421 -432 -420
rect -204 -421 -201 -418
rect -17 -420 -14 -401
rect 2 -410 5 -354
rect 32 -357 35 -349
rect 43 -349 46 -341
rect 43 -352 93 -349
rect 90 -356 93 -352
rect 107 -353 110 -322
rect 32 -360 83 -357
rect 80 -365 83 -360
rect 165 -365 168 -336
rect 80 -368 168 -365
rect 20 -397 26 -394
rect 2 -413 12 -410
rect 9 -420 12 -413
rect -435 -424 -434 -421
rect -204 -424 -162 -421
rect -17 -423 3 -420
rect 9 -423 32 -420
rect -165 -454 -162 -424
rect 0 -430 3 -423
rect 0 -433 19 -430
rect -544 -464 -541 -463
rect -567 -466 -541 -464
rect -570 -467 -541 -466
rect -506 -485 -503 -463
rect -471 -466 -441 -463
rect -384 -463 -347 -460
rect -235 -460 -198 -457
rect -235 -461 -232 -460
rect -258 -463 -232 -461
rect -384 -464 -381 -463
rect -407 -466 -381 -464
rect -410 -467 -381 -466
rect -506 -488 -473 -485
rect -346 -485 -343 -463
rect -261 -464 -232 -463
rect -197 -482 -194 -460
rect -83 -460 -46 -457
rect -83 -461 -80 -460
rect -106 -463 -80 -461
rect -109 -464 -80 -463
rect -346 -488 -313 -485
rect -197 -485 -164 -482
rect -131 -505 -128 -472
rect -45 -482 -42 -460
rect -45 -485 -12 -482
rect 29 -505 32 -423
rect -131 -508 32 -505
rect -139 -520 -132 -519
rect -139 -525 -138 -520
rect -133 -523 -79 -520
rect -133 -525 -132 -523
rect -139 -526 -132 -525
rect -82 -538 -79 -523
rect -539 -682 -536 -672
rect -120 -682 -117 -670
rect -614 -685 -540 -683
rect -618 -686 -540 -685
rect -535 -686 -458 -683
rect -453 -686 -374 -683
rect -369 -686 -292 -683
rect -287 -686 -206 -683
rect -201 -686 -121 -683
rect -116 -686 -38 -683
rect -33 -686 46 -683
<< m234contact >>
rect -91 -126 -86 -121
rect -294 -206 -289 -201
rect -227 -229 -222 -224
rect -294 -313 -289 -308
rect -398 -358 -393 -353
rect -387 -386 -382 -381
rect -18 -346 -13 -341
rect -420 -450 -415 -445
<< m4contact >>
rect -470 -330 -465 -325
rect -506 -335 -501 -330
rect -134 -252 -129 -247
rect -362 -342 -357 -337
rect -186 -413 -181 -408
rect 5 -359 10 -354
rect 106 -358 111 -353
rect 15 -398 20 -393
<< metal4 >>
rect -293 -308 -290 -206
rect -222 -229 -217 -225
rect -220 -235 -217 -229
rect -220 -238 -134 -235
rect -137 -252 -134 -238
rect -465 -328 -369 -325
rect -501 -334 -477 -331
rect -480 -354 -477 -334
rect -372 -339 -369 -328
rect -90 -334 -87 -126
rect -90 -337 -14 -334
rect -372 -342 -362 -339
rect -17 -341 -14 -337
rect -480 -357 -398 -354
rect 10 -358 106 -355
rect -386 -437 -383 -386
rect 7 -398 15 -395
rect 7 -405 10 -398
rect 7 -408 18 -405
rect -181 -412 -169 -409
rect -172 -417 -169 -412
rect 15 -417 18 -408
rect -172 -420 18 -417
rect -419 -440 -383 -437
rect -419 -445 -416 -440
<< m345contact >>
rect -215 -217 -210 -212
rect -136 -275 -131 -270
rect -36 -353 -31 -348
rect -434 -426 -429 -421
<< metal5 >>
rect -214 -230 -211 -217
rect -214 -233 -121 -230
rect -191 -243 -139 -240
rect -191 -314 -188 -243
rect -181 -250 -146 -247
rect -181 -311 -178 -250
rect -149 -280 -146 -250
rect -142 -270 -139 -243
rect -142 -274 -136 -270
rect -124 -280 -121 -233
rect -149 -283 -121 -280
rect -181 -314 -94 -311
rect -218 -317 -188 -314
rect -218 -360 -215 -317
rect -97 -349 -94 -314
rect -97 -352 -36 -349
rect -350 -363 -215 -360
rect -350 -422 -347 -363
rect -429 -425 -347 -422
<< labels >>
rlabel metal1 -547 -447 -547 -447 1 b0_inv
rlabel metal1 -444 -474 -438 -471 7 g0_inv
rlabel metal1 -478 -463 -474 -460 1 p0_inv
rlabel metal1 -541 -509 -539 -506 1 b0
rlabel metal2 -579 -449 -577 -447 3 mid_s0
rlabel metal1 -566 -468 -564 -466 1 a0
rlabel metal1 -499 -525 -499 -524 1 vdd
rlabel metal1 -489 -443 -489 -443 5 gnd
rlabel metal1 -569 -437 -569 -437 1 gnd
rlabel metal1 -600 -416 -598 -414 1 s0
rlabel metal1 -612 -417 -610 -415 1 c0
rlabel metal1 -579 -418 -576 -416 1 mid_s0
rlabel metal1 -444 -405 -438 -402 7 c1
rlabel metal1 -471 -405 -467 -403 1 g0_inv
rlabel metal1 -451 -434 -451 -434 1 gnd
rlabel metal1 -477 -398 -475 -395 1 temp100
rlabel metal1 -504 -420 -504 -420 1 gnd
rlabel metal1 -529 -376 -527 -373 1 c0_inv
rlabel metal1 -544 -377 -542 -375 3 c0
rlabel metal1 -354 -505 -354 -505 1 vdd
rlabel metal1 -329 -443 -329 -443 5 gnd
rlabel metal1 -339 -525 -339 -524 1 vdd
rlabel metal1 -300 -515 -300 -515 1 vdd
rlabel metal2 -419 -449 -417 -447 3 mid_s1
rlabel metal1 -406 -468 -404 -466 1 a1
rlabel metal1 -381 -509 -379 -506 1 b1
rlabel metal1 -318 -463 -314 -460 1 p1_inv
rlabel metal1 -284 -474 -278 -471 7 g1_inv
rlabel m2contact -380 -448 -378 -446 1 b1_inv
rlabel metal1 -406 -404 -404 -402 1 s1
rlabel metal1 -366 -366 -366 -366 5 vdd
rlabel metal1 -325 -268 -325 -267 5 vdd
rlabel metal1 -335 -349 -335 -349 1 gnd
rlabel metal1 -324 -326 -320 -324 7 p1_inv
rlabel metal1 -323 -332 -318 -330 7 p0_inv
rlabel metal1 -351 -328 -347 -326 3 temp101
rlabel metal1 -381 -274 -381 -274 5 vdd
rlabel metal1 -390 -347 -390 -347 1 gnd
rlabel metal1 -374 -318 -370 -317 1 c0
rlabel metal1 -418 -317 -416 -315 1 temp102
rlabel metal1 -407 -245 -407 -245 3 gnd
rlabel metal1 -326 -255 -325 -255 7 vdd
rlabel metal1 -385 -219 -382 -216 1 temp103
rlabel metal1 -298 -220 -298 -220 5 vdd
rlabel metal1 -289 -293 -289 -293 1 gnd
rlabel metal1 -306 -264 -306 -264 1 g1_inv
rlabel metal1 -282 -264 -276 -261 7 temp104
rlabel metal1 -260 -220 -260 -219 5 vdd
rlabel metal1 -250 -301 -250 -301 1 gnd
rlabel metal1 -223 -279 -221 -277 1 c2
rlabel metal1 -390 -263 -387 -260 1 g0_inv
rlabel metal1 -521 -403 -516 -400 1 p0_inv
rlabel metal1 -232 -506 -230 -503 1 b2
rlabel metal1 -257 -465 -255 -463 1 a2
rlabel metal2 -270 -446 -268 -444 3 mid_s2
rlabel m2contact -231 -445 -229 -443 1 b2_inv
rlabel metal1 -169 -460 -165 -457 1 p2_inv
rlabel metal1 -135 -471 -129 -468 7 g2_inv
rlabel metal1 -151 -512 -151 -512 1 vdd
rlabel metal1 -190 -522 -190 -521 1 vdd
rlabel metal1 -180 -440 -180 -440 5 gnd
rlabel metal1 -205 -502 -205 -502 1 vdd
rlabel metal1 -269 -352 -267 -350 1 s2
rlabel metal1 -238 -373 -238 -373 1 gnd
rlabel metal1 -104 -187 -104 -186 5 vdd
rlabel metal1 -94 -268 -94 -268 1 gnd
rlabel metal1 -48 -193 -48 -193 5 vdd
rlabel metal1 -39 -266 -39 -266 1 gnd
rlabel metal1 -22 -164 -22 -164 7 gnd
rlabel metal1 -104 -174 -103 -174 3 vdd
rlabel metal1 -131 -139 -131 -139 5 vdd
rlabel metal1 -140 -212 -140 -212 1 gnd
rlabel metal1 -169 -139 -169 -138 5 vdd
rlabel metal1 -179 -220 -179 -220 1 gnd
rlabel metal1 -208 -198 -206 -196 1 c3
rlabel metal1 -153 -183 -147 -180 1 temp108
rlabel metal1 -13 -236 -11 -234 1 temp106
rlabel metal1 -59 -237 -55 -236 1 c1
rlabel metal1 -82 -247 -78 -245 1 temp105
rlabel metal1 -109 -245 -105 -243 1 p2_inv
rlabel metal1 -47 -138 -44 -135 1 temp107
rlabel metal1 -124 -184 -122 -182 1 g2_inv
rlabel metal1 -41 -180 -38 -177 1 g1_inv
rlabel metal1 -107 -250 -107 -250 1 p1_inv
rlabel metal1 -118 -322 -118 -321 5 vdd
rlabel metal1 -128 -403 -128 -403 1 gnd
rlabel metal1 -117 -380 -113 -378 7 p3_inv
rlabel metal1 -143 -382 -142 -380 3 temp109
rlabel metal1 -160 -327 -160 -327 5 vdd
rlabel metal1 -169 -400 -169 -400 1 gnd
rlabel metal1 -153 -365 -150 -362 1 temp101
rlabel metal1 -197 -370 -195 -368 1 p4
rlabel metal1 -53 -502 -53 -502 1 vdd
rlabel metal1 -28 -440 -28 -440 5 gnd
rlabel metal1 -38 -522 -38 -521 1 vdd
rlabel metal1 1 -512 1 -512 1 vdd
rlabel m2contact -79 -445 -77 -443 1 b3_inv
rlabel metal2 -118 -446 -116 -444 3 mid_s3
rlabel metal1 -105 -465 -103 -463 1 a3
rlabel metal1 17 -471 23 -468 7 g3_inv
rlabel metal1 -17 -460 -13 -457 1 p3_inv
rlabel m123contact -114 -385 -114 -385 1 p2_inv
rlabel metal1 -240 -316 -240 -316 1 vdd
rlabel metal3 -34 -394 -34 -394 1 in2
rlabel metal1 -76 -415 -76 -415 1 gnd
rlabel metal1 -85 -356 -85 -356 5 vdd
rlabel metal1 -47 -394 -45 -392 1 s3
rlabel metal1 151 -390 153 -387 1 g4_inv
rlabel metal1 174 -374 174 -374 7 gnd
rlabel metal1 92 -364 93 -364 3 vdd
rlabel metal1 201 -329 207 -326 7 temp112
rlabel metal1 175 -330 177 -327 1 g3_inv
rlabel metal1 194 -358 194 -358 1 gnd
rlabel metal1 185 -285 185 -285 5 vdd
rlabel m2contact 117 -328 117 -328 1 p3_inv
rlabel metal1 158 -322 160 -320 1 temp111
rlabel metal1 131 -344 131 -344 1 gnd
rlabel metal1 121 -263 121 -262 5 vdd
rlabel metal1 2 -312 2 -312 1 temp110
rlabel metal1 42 -311 54 -308 1 temp104
rlabel metal1 48 -316 48 -316 1 temp109
rlabel metal1 41 -253 41 -252 5 vdd
rlabel metal1 31 -334 31 -334 1 gnd
rlabel metal1 96 -316 96 -314 1 temp110
rlabel metal1 69 -346 69 -346 1 gnd
rlabel metal1 60 -273 60 -273 5 vdd
rlabel metal1 55 -398 55 -398 5 vdd
rlabel metal1 64 -471 64 -471 1 gnd
rlabel metal1 46 -436 48 -433 3 p4
rlabel metal1 45 -443 48 -440 3 c0
rlabel metal1 89 -398 89 -398 5 vdd
rlabel metal1 98 -471 98 -471 1 gnd
rlabel metal1 81 -442 83 -441 1 temp113
rlabel m2contact 79 -436 82 -433 1 g4_inv
rlabel metal1 105 -442 111 -439 7 c4
rlabel m2contact -80 -507 -78 -504 1 b3
rlabel metal1 -472 -656 -472 -656 7 gnd
rlabel metal1 -551 -655 -551 -655 7 gnd
rlabel metal1 -616 -673 -616 -673 3 vdd
rlabel metal1 -390 -653 -390 -653 7 gnd
rlabel m2contact -383 -676 -383 -676 7 clk
rlabel metal1 -455 -671 -455 -671 3 vdd
rlabel metal1 -306 -654 -306 -654 7 gnd
rlabel m2contact -299 -677 -299 -677 7 clk
rlabel metal1 -371 -672 -371 -672 3 vdd
rlabel metal1 -224 -653 -224 -653 7 gnd
rlabel m2contact -217 -676 -217 -676 7 clk
rlabel metal1 -289 -671 -289 -671 3 vdd
rlabel metal1 -138 -653 -138 -653 7 gnd
rlabel m2contact -131 -676 -131 -676 7 clk
rlabel metal1 -203 -671 -203 -671 3 vdd
rlabel metal1 -53 -654 -53 -654 7 gnd
rlabel m2contact -46 -677 -46 -677 7 clk
rlabel metal1 -118 -672 -118 -672 3 vdd
rlabel metal1 30 -654 30 -654 7 gnd
rlabel m2contact 37 -677 37 -677 7 clk
rlabel metal1 114 -654 114 -654 7 gnd
rlabel m2contact 121 -677 121 -677 7 clk
rlabel metal1 49 -672 49 -672 3 vdd
rlabel metal1 -580 -680 -578 -678 1 c0_in
rlabel metal1 -501 -681 -499 -679 1 a0_in
rlabel metal1 -419 -678 -417 -676 1 b0_in
rlabel metal1 -335 -679 -333 -677 1 a1_in
rlabel metal1 -253 -678 -251 -676 1 b1_in
rlabel metal1 -167 -678 -165 -676 1 a2_in
rlabel metal1 -82 -679 -80 -677 1 b2_in
rlabel metal1 1 -679 3 -677 1 a3_in
rlabel metal1 85 -679 87 -677 1 b3_in
rlabel metal1 -35 -672 -35 -672 3 vdd
rlabel metal1 -537 -674 -537 -674 3 vdd
rlabel m2contact -464 -679 -464 -679 7 clk
rlabel m2contact -544 -676 -544 -676 7 clk
rlabel metal1 -631 -345 -631 -345 3 vdd
rlabel metal1 -559 -350 -559 -350 7 clk
rlabel metal1 -566 -327 -566 -327 7 gnd
rlabel m2contact -595 -352 -593 -349 1 s0
rlabel metal1 -593 -217 -593 -217 7 s0_out
rlabel metal1 -632 -204 -632 -204 3 vdd
rlabel metal1 -574 -203 -574 -203 7 gnd
rlabel metal1 -595 -193 -595 -193 7 s0_inv
rlabel metal1 -531 -307 -531 -307 3 vdd
rlabel metal1 -459 -312 -459 -312 7 clk
rlabel metal1 -466 -289 -466 -289 7 gnd
rlabel metal1 -532 -166 -532 -166 3 vdd
rlabel metal1 -474 -165 -474 -165 7 gnd
rlabel m2contact -495 -314 -493 -311 1 s1
rlabel metal1 -495 -156 -495 -156 1 s1_inv
rlabel metal1 -496 -180 -492 -178 1 s1_out
rlabel metal1 -272 -45 -272 -45 7 gnd
rlabel metal1 -330 -46 -330 -46 3 vdd
rlabel metal1 -264 -169 -264 -169 7 gnd
rlabel metal1 -257 -192 -257 -192 7 clk
rlabel metal1 -329 -187 -329 -187 3 vdd
rlabel metal1 -294 -61 -290 -58 1 s2_out
rlabel metal1 -294 -36 -292 -34 1 s2_inv
rlabel metal1 -69 43 -69 43 7 gnd
rlabel metal1 -127 42 -127 42 3 vdd
rlabel metal1 -61 -81 -61 -81 7 gnd
rlabel metal1 -54 -104 -54 -104 7 clk
rlabel metal1 -126 -99 -126 -99 3 vdd
rlabel metal1 -91 28 -87 30 1 s3_out
rlabel metal1 -90 52 -90 54 1 s3_inv
rlabel metal1 17 -230 17 -230 3 vdd
rlabel metal1 89 -235 89 -235 7 clk
rlabel metal1 82 -212 82 -212 7 gnd
rlabel metal1 16 -89 16 -89 3 vdd
rlabel metal1 74 -88 74 -88 7 gnd
rlabel metal1 53 -237 55 -232 1 c4
rlabel metal1 53 -103 55 -101 1 c4_out
rlabel metal1 52 -79 55 -77 1 c4_inv
<< end >>
