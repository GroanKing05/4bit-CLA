magic
tech scmos
timestamp 1731433869
<< nwell >>
rect -61 136 81 168
rect -61 46 81 78
<< ntransistor >>
rect -50 110 -48 130
rect -26 110 -24 130
rect 0 116 2 126
rect 18 110 20 130
rect 27 110 29 130
rect 43 110 45 130
rect 52 110 54 130
rect 68 116 70 126
rect -50 20 -48 40
rect -26 20 -24 40
rect 0 26 2 36
rect 18 20 20 40
rect 27 20 29 40
rect 43 20 45 40
rect 52 20 54 40
rect 68 26 70 36
<< ptransistor >>
rect -50 142 -48 162
rect -42 142 -40 162
rect -26 142 -24 162
rect -18 142 -16 162
rect 0 142 2 162
rect 18 142 20 162
rect 43 142 45 162
rect 68 142 70 162
rect -50 52 -48 72
rect -42 52 -40 72
rect -26 52 -24 72
rect -18 52 -16 72
rect 0 52 2 72
rect 18 52 20 72
rect 43 52 45 72
rect 68 52 70 72
<< ndiffusion >>
rect -55 114 -50 130
rect -51 110 -50 114
rect -48 126 -47 130
rect -48 110 -43 126
rect -31 114 -26 130
rect -27 110 -26 114
rect -24 126 -23 130
rect -24 110 -19 126
rect -5 120 0 126
rect -1 116 0 120
rect 2 122 3 126
rect 2 116 7 122
rect 13 114 18 130
rect 17 110 18 114
rect 20 110 27 130
rect 29 126 30 130
rect 29 110 34 126
rect 38 114 43 130
rect 42 110 43 114
rect 45 110 52 130
rect 54 126 55 130
rect 54 110 59 126
rect 63 120 68 126
rect 67 116 68 120
rect 70 122 71 126
rect 70 116 75 122
rect -55 24 -50 40
rect -51 20 -50 24
rect -48 36 -47 40
rect -48 20 -43 36
rect -31 24 -26 40
rect -27 20 -26 24
rect -24 36 -23 40
rect -24 20 -19 36
rect -5 30 0 36
rect -1 26 0 30
rect 2 32 3 36
rect 2 26 7 32
rect 13 24 18 40
rect 17 20 18 24
rect 20 20 27 40
rect 29 36 30 40
rect 29 20 34 36
rect 38 24 43 40
rect 42 20 43 24
rect 45 20 52 40
rect 54 36 55 40
rect 54 20 59 36
rect 63 30 68 36
rect 67 26 68 30
rect 70 32 71 36
rect 70 26 75 32
<< pdiffusion >>
rect -51 158 -50 162
rect -55 142 -50 158
rect -48 142 -42 162
rect -40 146 -35 162
rect -40 142 -39 146
rect -27 158 -26 162
rect -31 142 -26 158
rect -24 142 -18 162
rect -16 146 -11 162
rect -16 142 -15 146
rect -1 158 0 162
rect -5 142 0 158
rect 2 146 7 162
rect 2 142 3 146
rect 17 158 18 162
rect 13 142 18 158
rect 20 146 25 162
rect 20 142 21 146
rect 42 158 43 162
rect 38 142 43 158
rect 45 146 50 162
rect 45 142 46 146
rect 67 158 68 162
rect 63 142 68 158
rect 70 146 75 162
rect 70 142 71 146
rect -51 68 -50 72
rect -55 52 -50 68
rect -48 52 -42 72
rect -40 56 -35 72
rect -40 52 -39 56
rect -27 68 -26 72
rect -31 52 -26 68
rect -24 52 -18 72
rect -16 56 -11 72
rect -16 52 -15 56
rect -1 68 0 72
rect -5 52 0 68
rect 2 56 7 72
rect 2 52 3 56
rect 17 68 18 72
rect 13 52 18 68
rect 20 56 25 72
rect 20 52 21 56
rect 42 68 43 72
rect 38 52 43 68
rect 45 56 50 72
rect 45 52 46 56
rect 67 68 68 72
rect 63 52 68 68
rect 70 56 75 72
rect 70 52 71 56
<< ndcontact >>
rect -55 110 -51 114
rect -47 126 -43 130
rect -31 110 -27 114
rect -23 126 -19 130
rect -5 116 -1 120
rect 3 122 7 126
rect 13 110 17 114
rect 30 126 34 130
rect 38 110 42 114
rect 55 126 59 130
rect 63 116 67 120
rect 71 122 75 126
rect -55 20 -51 24
rect -47 36 -43 40
rect -31 20 -27 24
rect -23 36 -19 40
rect -5 26 -1 30
rect 3 32 7 36
rect 13 20 17 24
rect 30 36 34 40
rect 38 20 42 24
rect 55 36 59 40
rect 63 26 67 30
rect 71 32 75 36
<< pdcontact >>
rect -55 158 -51 162
rect -39 142 -35 146
rect -31 158 -27 162
rect -15 142 -11 146
rect -5 158 -1 162
rect 3 142 7 146
rect 13 158 17 162
rect 21 142 25 146
rect 38 158 42 162
rect 46 142 50 146
rect 63 158 67 162
rect 71 142 75 146
rect -55 68 -51 72
rect -39 52 -35 56
rect -31 68 -27 72
rect -15 52 -11 56
rect -5 68 -1 72
rect 3 52 7 56
rect 13 68 17 72
rect 21 52 25 56
rect 38 68 42 72
rect 46 52 50 56
rect 63 68 67 72
rect 71 52 75 56
<< polysilicon >>
rect -50 162 -48 166
rect -42 162 -40 166
rect -26 162 -24 166
rect -18 162 -16 166
rect 0 162 2 166
rect 18 162 20 165
rect 43 162 45 165
rect 68 162 70 166
rect -50 130 -48 142
rect -50 107 -48 110
rect -42 101 -40 142
rect -26 130 -24 142
rect -26 107 -24 110
rect -41 98 -40 101
rect -18 98 -16 142
rect 0 126 2 142
rect 18 130 20 142
rect 27 130 29 134
rect 43 130 45 142
rect 52 130 54 134
rect 0 112 2 116
rect 68 126 70 142
rect 68 112 70 116
rect 18 105 20 110
rect 27 96 29 110
rect 43 105 45 110
rect 52 96 54 110
rect -50 72 -48 76
rect -42 72 -40 76
rect -26 72 -24 76
rect -18 72 -16 76
rect 0 72 2 76
rect 18 72 20 75
rect 43 72 45 75
rect 68 72 70 76
rect -50 40 -48 52
rect -50 17 -48 20
rect -42 11 -40 52
rect -26 40 -24 52
rect -26 17 -24 20
rect -41 8 -40 11
rect -18 8 -16 52
rect 0 36 2 52
rect 18 40 20 52
rect 27 40 29 44
rect 43 40 45 52
rect 52 40 54 44
rect 0 22 2 26
rect 68 36 70 52
rect 68 22 70 26
rect 18 15 20 20
rect 27 6 29 20
rect 43 15 45 20
rect 52 6 54 20
<< polycontact >>
rect -54 131 -50 135
rect -30 131 -26 135
rect -45 97 -41 101
rect -22 97 -18 101
rect -4 130 0 134
rect 14 131 18 135
rect 39 131 43 135
rect 64 130 68 134
rect 23 97 27 101
rect 48 97 52 101
rect -54 41 -50 45
rect -30 41 -26 45
rect -45 7 -41 11
rect -22 7 -18 11
rect -4 40 0 44
rect 14 41 18 45
rect 39 41 43 45
rect 64 40 68 44
rect 23 7 27 11
rect 48 7 52 11
<< metal1 >>
rect -55 169 78 172
rect -55 162 -52 169
rect -31 162 -28 169
rect -5 162 -2 169
rect 13 162 16 169
rect 38 162 41 169
rect 63 162 66 169
rect -61 131 -54 134
rect -38 134 -35 142
rect -46 131 -30 134
rect -14 134 -11 142
rect 25 142 34 145
rect 50 142 59 145
rect 3 134 7 142
rect -22 131 -4 134
rect -46 130 -43 131
rect -22 130 -19 131
rect 3 131 14 134
rect 31 134 34 142
rect 31 131 39 134
rect 56 134 59 142
rect 71 134 75 142
rect 56 131 64 134
rect 3 126 7 131
rect 31 130 34 131
rect 56 130 59 131
rect 71 131 78 134
rect 71 126 75 131
rect -55 107 -52 110
rect -31 107 -28 110
rect -5 107 -2 116
rect 13 107 16 110
rect 38 107 41 110
rect 63 107 66 116
rect -55 104 66 107
rect -61 97 -45 100
rect -41 97 -22 100
rect -18 97 23 100
rect 27 97 48 100
rect -55 79 78 82
rect -55 72 -52 79
rect -31 72 -28 79
rect -5 72 -2 79
rect 13 72 16 79
rect 38 72 41 79
rect 63 72 66 79
rect -61 41 -54 44
rect -38 44 -35 52
rect -46 41 -30 44
rect -14 44 -11 52
rect 25 52 34 55
rect 50 52 59 55
rect 3 44 7 52
rect -22 41 -4 44
rect -46 40 -43 41
rect -22 40 -19 41
rect 3 41 14 44
rect 31 44 34 52
rect 31 41 39 44
rect 56 44 59 52
rect 71 44 75 52
rect 56 41 64 44
rect 3 36 7 41
rect 31 40 34 41
rect 56 40 59 41
rect 71 41 78 44
rect 71 36 75 41
rect -55 17 -52 20
rect -31 17 -28 20
rect -5 17 -2 26
rect 13 17 16 20
rect 38 17 41 20
rect 63 17 66 26
rect -55 14 66 17
rect -61 7 -45 10
rect -41 7 -22 10
rect -18 7 23 10
rect 27 7 48 10
<< labels >>
rlabel metal1 -54 170 -54 170 5 vdd
rlabel metal1 -59 98 -59 98 1 clk
rlabel metal1 -36 105 -36 105 1 gnd
rlabel metal1 -54 80 -54 80 5 vdd
rlabel metal1 -59 8 -59 8 1 clk
rlabel metal1 -36 15 -36 15 1 gnd
rlabel metal1 -60 132 -58 134 3 a0_in
rlabel metal1 73 131 77 134 1 a0
rlabel metal1 -61 42 -56 44 3 b0_in
rlabel metal1 74 41 77 44 1 b0
<< end >>
