magic
tech scmos
timestamp 1731391111
<< nwell >>
rect -60 18 -28 43
rect -21 23 12 55
<< ntransistor >>
rect -76 30 -66 32
rect -10 6 -8 16
rect -1 6 1 16
<< ptransistor >>
rect -54 30 -34 32
rect -10 29 -8 49
rect -1 29 1 49
<< ndiffusion >>
rect -72 33 -66 37
rect -76 32 -66 33
rect -76 29 -66 30
rect -76 25 -70 29
rect -15 10 -10 16
rect -11 6 -10 10
rect -8 12 -7 16
rect -3 12 -1 16
rect -8 6 -1 12
rect 1 12 2 16
rect 1 6 6 12
<< pdiffusion >>
rect -11 45 -10 49
rect -54 33 -38 37
rect -54 32 -34 33
rect -54 29 -34 30
rect -15 29 -10 45
rect -8 35 -1 49
rect -8 31 -7 35
rect -3 31 -1 35
rect -8 29 -1 31
rect 1 33 6 49
rect 1 29 2 33
rect -50 25 -34 29
<< ndcontact >>
rect -76 33 -72 37
rect -70 25 -66 29
rect -15 6 -11 10
rect -7 12 -3 16
rect 2 12 6 16
<< pdcontact >>
rect -15 45 -11 49
rect -38 33 -34 37
rect -7 31 -3 35
rect 2 29 6 33
rect -54 25 -50 29
<< polysilicon >>
rect -10 49 -8 52
rect -1 49 1 61
rect -80 30 -76 32
rect -66 30 -54 32
rect -34 30 -30 32
rect -10 16 -8 29
rect -1 23 1 29
rect -1 16 1 20
rect -10 3 -8 6
rect -1 4 1 6
rect 0 0 1 4
rect -1 -1 1 0
<< polycontact >>
rect -5 56 -1 60
rect -65 32 -61 36
rect -14 18 -10 22
rect -4 0 0 4
<< metal1 >>
rect -27 56 -5 59
rect -27 49 -24 56
rect -64 46 -15 49
rect -84 34 -76 37
rect -64 36 -61 46
rect -34 34 -24 37
rect -66 25 -54 28
rect -6 28 -3 31
rect -64 17 -61 25
rect -20 18 -14 21
rect -64 14 -31 17
rect -6 16 -3 23
rect -34 11 -31 14
rect 2 22 5 29
rect 2 20 12 22
rect 2 19 9 20
rect 2 16 5 19
rect -34 9 -18 11
rect -34 8 -15 9
rect -21 6 -15 8
rect -21 3 -18 6
rect -21 0 -4 3
<< m2contact >>
rect -7 23 -2 28
<< metal2 >>
rect -2 24 14 27
<< m123contact >>
rect -25 17 -20 22
rect 9 15 14 20
<< metal3 >>
rect -20 20 12 21
rect -20 18 9 20
<< labels >>
rlabel metal1 -63 26 -63 26 3 in1_inv
rlabel metal1 -64 39 -62 42 5 in1
rlabel metal1 -83 36 -83 36 3 gnd
rlabel metal1 -26 36 -26 36 1 vdd
rlabel metal1 -5 22 -5 22 1 out
rlabel metal3 7 21 7 21 1 in2
<< end >>
