* SPICE3 file created from bit1gen.ext - technology: scmos
* Adds 1 bit and generates s0 and c1
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global gnd vdd

M1000 vdd mid_s0 a_6_n255# w_22_n262# CMOSP w=20 l=2
+  ad=1240 pd=584 as=100 ps=50
M1001 vdd g0_inv c1 w_37_n150# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1002 a_123_n204# temp100 gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=600 ps=340
M1003 s0 c0 mid_s0 w_61_n257# CMOSP w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1004 g0_inv b0 vdd w_n37_n170# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1005 temp100 a_74_n192# vdd w_37_n150# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 gnd a0 a_n24_n202# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1007 gnd b0 a_n84_n281# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1008 gnd mid_s0 a_6_n255# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1009 c0 mid_s0 s0 w_61_n257# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 a_n84_n281# a0 mid_s0 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1011 temp100 a_74_n192# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1012 mid_s0 a_n84_n281# a0 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1013 c1 temp100 vdd w_37_n150# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 vdd a0 g0_inv w_n37_n170# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 b0 a0 mid_s0 w_n95_n257# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1016 a_10_n164# b0 vdd w_n37_n170# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1017 c0_inv c0 vdd w_37_n150# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1018 p0_inv b0 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1019 mid_s0 b0 a0 w_n95_n257# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1020 vdd b0 a_n84_n281# w_n55_n262# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1021 c0_inv c0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1022 p0_inv a0 a_10_n164# w_n37_n170# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1023 gnd a0 p0_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 a_74_n192# c0_inv a_74_n164# w_37_n150# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1025 gnd c0_inv a_74_n192# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1026 c1 g0_inv a_123_n204# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1027 a_n24_n202# b0 g0_inv Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1028 s0 c0 a_6_n255# Gnd CMOSN w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1029 a_74_n164# p0_inv vdd w_37_n150# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 a_74_n192# p0_inv gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 c0 a_6_n255# s0 Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 c0 c0_inv 0.04fF
C1 gnd a_6_n255# 0.02fF
C2 w_n37_n170# g0_inv 0.30fF
C3 b0 p0_inv 0.02fF
C4 g0_inv c1 0.10fF
C5 w_n37_n170# p0_inv 0.02fF
C6 w_n55_n262# b0 0.07fF
C7 w_n95_n257# a0 0.24fF
C8 w_37_n150# c0 0.07fF
C9 g0_inv a_74_n164# 0.01fF
C10 g0_inv a_10_n164# 0.01fF
C11 vdd gnd 0.42fF
C12 w_n37_n170# b0 0.14fF
C13 w_22_n262# a_6_n255# 0.02fF
C14 b0 mid_s0 0.25fF
C15 c0_inv gnd 0.03fF
C16 mid_s0 s0 0.00fF
C17 c0 g0_inv 0.07fF
C18 a0 vdd 0.12fF
C19 w_37_n150# temp100 0.09fF
C20 w_22_n262# vdd 0.11fF
C21 w_37_n150# vdd 0.14fF
C22 c0 p0_inv 0.12fF
C23 a_74_n192# temp100 0.04fF
C24 w_37_n150# c0_inv 0.12fF
C25 gnd a_74_n192# 0.04fF
C26 g0_inv temp100 0.31fF
C27 c0 s0 0.35fF
C28 w_n95_n257# b0 0.10fF
C29 g0_inv gnd 0.01fF
C30 w_61_n257# s0 0.17fF
C31 a0 a_n84_n281# 0.10fF
C32 c0 mid_s0 0.27fF
C33 vdd g0_inv 0.08fF
C34 w_61_n257# mid_s0 0.10fF
C35 c0_inv a_74_n192# 0.17fF
C36 w_n95_n257# mid_s0 0.18fF
C37 p0_inv gnd 0.16fF
C38 c0_inv g0_inv 0.12fF
C39 mid_s0 a_6_n255# 0.06fF
C40 b0 gnd 0.05fF
C41 a0 g0_inv 0.38fF
C42 b0 vdd 0.19fF
C43 w_37_n150# a_74_n192# 0.09fF
C44 w_n55_n262# vdd 0.11fF
C45 p0_inv c0_inv 0.25fF
C46 w_37_n150# g0_inv 0.39fF
C47 w_n37_n170# vdd 0.12fF
C48 a0 p0_inv 0.17fF
C49 gnd mid_s0 0.22fF
C50 vdd mid_s0 0.12fF
C51 b0 a0 0.71fF
C52 w_61_n257# c0 0.24fF
C53 w_37_n150# p0_inv 0.06fF
C54 g0_inv a_74_n192# 0.05fF
C55 c0 a_6_n255# 0.10fF
C56 w_n37_n170# a0 0.44fF
C57 a0 mid_s0 0.40fF
C58 b0 a_n84_n281# 0.06fF
C59 p0_inv a_74_n192# 0.02fF
C60 b0 a_n24_n202# 0.01fF
C61 w_22_n262# mid_s0 0.07fF
C62 w_n55_n262# a_n84_n281# 0.02fF
C63 c0 gnd 0.67fF
C64 p0_inv g0_inv 0.05fF
C65 w_37_n150# c1 0.04fF
C66 b0 g0_inv 0.26fF
C67 s0 Gnd 0.43fF
C68 a_6_n255# Gnd 0.38fF
C69 a_n84_n281# Gnd 0.38fF
C70 mid_s0 Gnd 1.09fF
C71 c1 Gnd 0.05fF
C72 temp100 Gnd 0.00fF
C73 a_74_n192# Gnd 0.18fF
C74 gnd Gnd 1.58fF
C75 g0_inv Gnd 1.03fF
C76 vdd Gnd 2.11fF
C77 c0_inv Gnd 0.09fF
C78 p0_inv Gnd 0.68fF
C79 c0 Gnd 0.24fF
C80 a0 Gnd 1.78fF
C81 b0 Gnd 1.19fF
C82 w_61_n257# Gnd 1.06fF
C83 w_22_n262# Gnd 0.84fF
C84 w_n55_n262# Gnd 0.84fF
C85 w_n95_n257# Gnd 1.06fF
C86 w_37_n150# Gnd 1.14fF
C87 w_n37_n170# Gnd 1.09fF

Vdd vdd gnd 'SUPPLY'
Va0 a0 gnd 1.8
Vb0 b0 gnd 1.8
Vc0 c0 gnd 1.8

.tran 100ps 400ns

.control
set hcopypscolor = 0
set color0=white 
set color1=black 

run

set curplottitle="2023112005_1_bit_adder"

plot a0, b0+2, c0+4, s0+6, c1+8
.endc