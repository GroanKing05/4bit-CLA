* SPICE3 file created from XOR2.ext - technology: scmos

.option scale=0.09u

M1000 out in2 in1 w_n191_n85# pfet w=20 l=2
+  ad=140 pd=54 as=100 ps=50
M1001 in2 in1 out w_n191_n85# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1002 gnd in1 in1_inv Gnd nfet w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1003 vdd in1 in1_inv w_n191_n85# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1004 in2 in1_inv out Gnd nfet w=10 l=2
+  ad=50 pd=30 as=70 ps=34
M1005 out in2 in1_inv Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in1 gnd 0.02fF
C1 in1 in2 0.07fF
C2 w_n191_n85# out 0.17fF
C3 w_n191_n85# in1_inv 0.02fF
C4 in1 out 0.00fF
C5 in1 in1_inv 0.06fF
C6 w_n191_n85# vdd 0.02fF
C7 w_n191_n85# in1 0.27fF
C8 in1_inv gnd 0.18fF
C9 in2 out 0.34fF
C10 in1 vdd 0.05fF
C11 in2 in1_inv 0.05fF
C12 w_n191_n85# in2 0.09fF
C13 gnd Gnd 0.06fF
C14 out Gnd 0.05fF
C15 vdd Gnd 0.04fF
C16 in1_inv Gnd 0.04fF
C17 in2 Gnd 0.24fF
C18 in1 Gnd 0.25fF
C19 w_n191_n85# Gnd 1.96fF
