magic
tech scmos
timestamp 1731591089
<< nwell >>
rect -20 -64 38 -42
rect -20 -74 87 -64
rect -91 -115 -30 -83
rect 4 -94 87 -74
rect 32 -96 87 -94
rect -45 -171 16 -170
rect -45 -182 53 -171
rect -45 -202 87 -182
rect 19 -214 87 -202
rect 19 -223 53 -214
<< ntransistor >>
rect -9 -90 -7 -80
rect 15 -116 17 -106
rect 25 -116 27 -106
rect 43 -112 45 -102
rect -80 -132 -78 -122
rect -71 -132 -69 -122
rect -43 -131 -41 -121
rect 64 -128 66 -108
rect 74 -128 76 -108
rect -34 -163 -32 -153
rect -25 -163 -23 -153
rect 3 -164 5 -154
rect 30 -159 32 -149
rect 40 -159 42 -149
rect 64 -170 66 -150
rect 74 -170 76 -150
<< ptransistor >>
rect -9 -68 -7 -48
rect -80 -109 -78 -89
rect -71 -109 -69 -89
rect -43 -109 -41 -89
rect 15 -88 17 -48
rect 25 -88 27 -48
rect 43 -90 45 -70
rect 64 -90 66 -70
rect 74 -90 76 -70
rect -34 -196 -32 -176
rect -25 -196 -23 -176
rect 3 -196 5 -176
rect 30 -217 32 -177
rect 40 -217 42 -177
rect 64 -208 66 -188
rect 74 -208 76 -188
<< ndiffusion >>
rect -14 -86 -9 -80
rect -10 -90 -9 -86
rect -7 -84 -6 -80
rect -7 -90 -2 -84
rect 10 -112 15 -106
rect 14 -116 15 -112
rect 17 -110 19 -106
rect 23 -110 25 -106
rect 17 -116 25 -110
rect 27 -112 32 -106
rect 38 -108 43 -102
rect 42 -112 43 -108
rect 45 -106 46 -102
rect 45 -112 50 -106
rect 27 -116 28 -112
rect -81 -126 -80 -122
rect -85 -132 -80 -126
rect -78 -126 -76 -122
rect -72 -126 -71 -122
rect -78 -132 -71 -126
rect -69 -128 -64 -122
rect -69 -132 -68 -128
rect -48 -127 -43 -121
rect -44 -131 -43 -127
rect -41 -127 -36 -121
rect -41 -131 -40 -127
rect 59 -124 64 -108
rect 63 -128 64 -124
rect 66 -128 74 -108
rect 76 -112 77 -108
rect 76 -128 81 -112
rect -39 -159 -34 -153
rect -35 -163 -34 -159
rect -32 -159 -25 -153
rect -32 -163 -30 -159
rect -26 -163 -25 -159
rect -23 -157 -22 -153
rect 29 -153 30 -149
rect -23 -163 -18 -157
rect 2 -158 3 -154
rect -2 -164 3 -158
rect 5 -158 6 -154
rect 5 -164 10 -158
rect 25 -159 30 -153
rect 32 -155 40 -149
rect 32 -159 34 -155
rect 38 -159 40 -155
rect 42 -153 43 -149
rect 42 -159 47 -153
rect 63 -154 64 -150
rect 59 -170 64 -154
rect 66 -170 74 -150
rect 76 -166 81 -150
rect 76 -170 77 -166
<< pdiffusion >>
rect -10 -52 -9 -48
rect -14 -68 -9 -52
rect -7 -64 -2 -48
rect -7 -68 -6 -64
rect 14 -52 15 -48
rect -85 -105 -80 -89
rect -81 -109 -80 -105
rect -78 -103 -71 -89
rect -78 -107 -76 -103
rect -72 -107 -71 -103
rect -78 -109 -71 -107
rect -69 -93 -68 -89
rect -69 -109 -64 -93
rect -44 -93 -43 -89
rect -48 -109 -43 -93
rect -41 -105 -36 -89
rect 10 -88 15 -52
rect 17 -88 25 -48
rect 27 -84 32 -48
rect 27 -88 28 -84
rect 42 -74 43 -70
rect -41 -109 -40 -105
rect 38 -90 43 -74
rect 45 -86 50 -70
rect 45 -90 46 -86
rect 63 -74 64 -70
rect 59 -90 64 -74
rect 66 -86 74 -70
rect 66 -90 68 -86
rect 72 -90 74 -86
rect 76 -74 77 -70
rect 76 -90 81 -74
rect -35 -180 -34 -176
rect -39 -196 -34 -180
rect -32 -178 -25 -176
rect -32 -182 -30 -178
rect -26 -182 -25 -178
rect -32 -196 -25 -182
rect -23 -192 -18 -176
rect -23 -196 -22 -192
rect -2 -192 3 -176
rect 2 -196 3 -192
rect 5 -180 6 -176
rect 5 -196 10 -180
rect 25 -213 30 -177
rect 29 -217 30 -213
rect 32 -217 40 -177
rect 42 -181 43 -177
rect 42 -217 47 -181
rect 59 -204 64 -188
rect 63 -208 64 -204
rect 66 -192 68 -188
rect 72 -192 74 -188
rect 66 -208 74 -192
rect 76 -204 81 -188
rect 76 -208 77 -204
<< ndcontact >>
rect -14 -90 -10 -86
rect -6 -84 -2 -80
rect 10 -116 14 -112
rect 19 -110 23 -106
rect 38 -112 42 -108
rect 46 -106 50 -102
rect 28 -116 32 -112
rect -85 -126 -81 -122
rect -76 -126 -72 -122
rect -68 -132 -64 -128
rect -48 -131 -44 -127
rect -40 -131 -36 -127
rect 59 -128 63 -124
rect 77 -112 81 -108
rect -39 -163 -35 -159
rect -30 -163 -26 -159
rect -22 -157 -18 -153
rect 25 -153 29 -149
rect -2 -158 2 -154
rect 6 -158 10 -154
rect 34 -159 38 -155
rect 43 -153 47 -149
rect 59 -154 63 -150
rect 77 -170 81 -166
<< pdcontact >>
rect -14 -52 -10 -48
rect -6 -68 -2 -64
rect 10 -52 14 -48
rect -85 -109 -81 -105
rect -76 -107 -72 -103
rect -68 -93 -64 -89
rect -48 -93 -44 -89
rect 28 -88 32 -84
rect 38 -74 42 -70
rect -40 -109 -36 -105
rect 46 -90 50 -86
rect 59 -74 63 -70
rect 68 -90 72 -86
rect 77 -74 81 -70
rect -39 -180 -35 -176
rect -30 -182 -26 -178
rect -22 -196 -18 -192
rect -2 -196 2 -192
rect 6 -180 10 -176
rect 25 -217 29 -213
rect 43 -181 47 -177
rect 59 -208 63 -204
rect 68 -192 72 -188
rect 77 -208 81 -204
<< polysilicon >>
rect -9 -48 -7 -44
rect 15 -48 17 -45
rect 25 -48 27 -45
rect -80 -89 -78 -77
rect -9 -80 -7 -68
rect -71 -89 -69 -86
rect -43 -89 -41 -85
rect 43 -70 45 -67
rect 64 -70 66 -66
rect 74 -70 76 -66
rect -9 -94 -7 -90
rect 15 -106 17 -88
rect 25 -106 27 -88
rect 43 -102 45 -90
rect -80 -115 -78 -109
rect -80 -122 -78 -118
rect -71 -122 -69 -109
rect -43 -121 -41 -109
rect 64 -108 66 -90
rect 74 -108 76 -90
rect 43 -115 45 -112
rect 15 -119 17 -116
rect 25 -119 27 -116
rect -80 -134 -78 -132
rect -80 -138 -79 -134
rect -71 -135 -69 -132
rect -43 -135 -41 -131
rect 64 -132 66 -128
rect 74 -132 76 -128
rect -80 -139 -78 -138
rect -34 -147 -32 -146
rect -34 -151 -33 -147
rect 30 -149 32 -146
rect 40 -149 42 -146
rect -34 -153 -32 -151
rect -25 -153 -23 -150
rect 3 -154 5 -150
rect -34 -167 -32 -163
rect -34 -176 -32 -170
rect -25 -176 -23 -163
rect 64 -150 66 -146
rect 74 -150 76 -146
rect 3 -176 5 -164
rect 30 -177 32 -159
rect 40 -177 42 -159
rect -34 -208 -32 -196
rect -25 -199 -23 -196
rect 3 -200 5 -196
rect 64 -188 66 -170
rect 74 -188 76 -170
rect 64 -212 66 -208
rect 74 -212 76 -208
rect 30 -220 32 -217
rect 40 -220 42 -217
<< polycontact >>
rect -78 -82 -74 -78
rect -13 -79 -9 -75
rect 11 -105 15 -101
rect 21 -99 25 -95
rect 39 -101 43 -97
rect 60 -101 64 -97
rect -69 -120 -65 -116
rect -47 -120 -43 -116
rect 70 -107 74 -103
rect -79 -138 -75 -134
rect -33 -151 -29 -147
rect 26 -164 30 -160
rect -23 -169 -19 -165
rect -1 -169 3 -165
rect 36 -170 40 -166
rect -32 -207 -28 -203
rect 60 -181 64 -177
rect 70 -175 74 -171
<< metal1 >>
rect -30 -41 41 -38
rect -30 -42 -20 -41
rect -30 -69 -26 -42
rect -14 -48 -11 -41
rect 10 -48 13 -41
rect 38 -60 41 -41
rect 38 -63 87 -60
rect -103 -73 -26 -69
rect -103 -146 -99 -73
rect -74 -82 -59 -79
rect -62 -89 -59 -82
rect -48 -89 -44 -73
rect -5 -75 -2 -68
rect 38 -70 41 -63
rect 59 -70 62 -63
rect 77 -70 81 -63
rect -17 -78 -13 -75
rect -5 -78 6 -75
rect -5 -80 -2 -78
rect -64 -92 -51 -89
rect -84 -116 -81 -109
rect -76 -110 -73 -107
rect -93 -118 -81 -116
rect -88 -119 -81 -118
rect -84 -122 -81 -119
rect -76 -122 -73 -115
rect -54 -116 -51 -92
rect -65 -120 -62 -117
rect -54 -119 -47 -116
rect -64 -133 -58 -129
rect -64 -135 -63 -133
rect -75 -138 -63 -135
rect -103 -150 -61 -146
rect -54 -147 -51 -119
rect -39 -125 -36 -109
rect -39 -127 -35 -125
rect -36 -130 -35 -127
rect -48 -136 -45 -131
rect -14 -136 -11 -90
rect 3 -95 6 -78
rect 3 -98 21 -95
rect 29 -97 32 -88
rect 47 -97 50 -90
rect 69 -91 72 -90
rect 69 -94 81 -91
rect 29 -100 39 -97
rect 8 -104 11 -101
rect 29 -102 32 -100
rect 47 -100 60 -97
rect 47 -102 50 -100
rect 20 -105 32 -102
rect 20 -106 23 -105
rect 78 -103 81 -94
rect 58 -107 70 -104
rect 78 -106 87 -103
rect 78 -108 81 -106
rect 10 -120 13 -116
rect 29 -120 32 -116
rect 38 -119 41 -112
rect -1 -123 37 -120
rect -1 -136 2 -123
rect 59 -132 62 -128
rect -48 -139 2 -136
rect 63 -136 84 -133
rect -2 -142 2 -139
rect -2 -145 62 -142
rect -65 -223 -61 -150
rect -29 -150 -17 -147
rect -18 -152 -17 -150
rect -18 -156 -12 -152
rect -2 -154 1 -145
rect 25 -149 28 -145
rect 44 -149 47 -145
rect 8 -154 11 -152
rect 10 -158 11 -154
rect 59 -150 62 -145
rect -50 -167 -47 -166
rect -38 -166 -35 -163
rect -42 -167 -35 -166
rect -50 -169 -35 -167
rect -50 -212 -47 -169
rect -38 -176 -35 -169
rect -30 -170 -27 -163
rect -19 -168 -16 -165
rect -8 -169 -1 -166
rect -8 -173 -5 -169
rect -30 -178 -27 -175
rect 7 -176 10 -158
rect 35 -160 38 -159
rect 23 -164 26 -161
rect 35 -161 47 -160
rect 35 -163 50 -161
rect 44 -164 55 -163
rect 19 -170 36 -167
rect 19 -173 22 -170
rect -8 -193 -5 -178
rect 44 -177 47 -164
rect 57 -174 70 -171
rect 78 -172 81 -170
rect 84 -172 87 -169
rect 78 -175 87 -172
rect 53 -181 60 -178
rect 53 -185 56 -181
rect 78 -184 81 -175
rect 69 -187 81 -184
rect 69 -188 72 -187
rect -18 -196 -5 -193
rect -16 -203 -13 -196
rect -28 -206 -13 -203
rect -2 -205 2 -196
rect -17 -212 -14 -206
rect -2 -208 22 -205
rect 19 -223 22 -208
rect -65 -224 22 -223
rect 59 -215 62 -208
rect 77 -215 81 -208
rect 25 -224 28 -217
rect 49 -218 87 -215
rect 49 -224 53 -218
rect -65 -227 53 -224
<< m2contact >>
rect -77 -115 -72 -110
rect -63 -138 -58 -133
rect -35 -130 -30 -125
rect 3 -106 8 -101
rect 37 -124 42 -119
rect 58 -137 63 -132
rect -55 -152 -50 -147
rect -17 -152 -12 -147
rect 11 -155 16 -150
rect -31 -175 -26 -170
rect -9 -178 -4 -173
rect 50 -163 55 -158
rect 18 -178 23 -173
rect 52 -175 57 -170
<< metal2 >>
rect -96 -111 -93 370
rect -96 -114 -77 -111
rect -61 -140 -58 -138
rect -34 -140 -31 -130
rect -61 -143 -31 -140
rect 3 -140 6 -106
rect 42 -123 58 -120
rect 55 -136 58 -123
rect 3 -143 54 -140
rect -12 -152 11 -151
rect -54 -171 -51 -152
rect -16 -154 11 -152
rect 51 -158 54 -143
rect -54 -174 -31 -171
rect 19 -171 22 -169
rect 19 -173 52 -171
rect -4 -177 18 -174
rect 23 -174 52 -173
<< m123contact >>
rect -22 -79 -17 -74
rect -93 -123 -88 -118
rect -62 -121 -57 -116
rect 53 -109 58 -104
rect -47 -167 -42 -162
rect 18 -164 23 -159
rect -16 -169 -11 -164
rect 84 -169 89 -164
rect 52 -190 57 -185
<< metal3 >>
rect -61 -78 -22 -75
rect -61 -116 -58 -78
rect -91 -118 -62 -117
rect -88 -120 -62 -118
rect -19 -164 18 -161
rect 54 -164 57 -109
rect -19 -165 -16 -164
rect -42 -167 -16 -165
rect -45 -168 -16 -167
rect 19 -186 22 -164
rect 54 -167 84 -164
rect 19 -189 52 -186
<< labels >>
rlabel metal1 -22 -148 -22 -148 1 b0_inv
rlabel metal1 81 -175 87 -172 7 g0_inv
rlabel metal1 47 -164 51 -161 1 p0_inv
rlabel metal1 -16 -210 -14 -207 1 b0
rlabel metal2 -54 -150 -52 -148 3 mid_s0
rlabel metal1 -41 -169 -39 -167 1 a0
rlabel metal1 26 -226 26 -225 1 vdd
rlabel metal1 36 -144 36 -144 5 gnd
rlabel metal1 -44 -138 -44 -138 1 gnd
rlabel metal1 -75 -117 -73 -115 1 s0
rlabel metal1 -87 -118 -85 -116 1 c0
rlabel metal1 -54 -119 -51 -117 1 mid_s0
rlabel metal1 81 -106 87 -103 7 c1
rlabel metal1 54 -106 58 -104 1 g0_inv
rlabel metal1 74 -135 74 -135 1 gnd
rlabel m2contact 4 -103 8 -102 1 p0_inv
rlabel metal1 48 -99 50 -96 1 temp100
rlabel metal1 21 -121 21 -121 1 gnd
rlabel metal1 -4 -77 -2 -74 1 c0_inv
rlabel metal1 -19 -78 -17 -76 3 c0
<< end >>
