magic
tech scmos
timestamp 1731424967
<< nwell >>
rect -72 77 -38 82
rect -72 71 -1 77
rect -72 45 21 71
rect -72 30 -38 45
rect -4 39 21 45
<< ntransistor >>
rect -61 8 -59 18
rect -51 8 -49 18
rect -24 13 -22 33
rect -14 13 -12 33
rect 7 23 9 33
<< ptransistor >>
rect -61 36 -59 76
rect -51 36 -49 76
rect -24 51 -22 71
rect -14 51 -12 71
rect 7 45 9 65
<< ndiffusion >>
rect -66 12 -61 18
rect -62 8 -61 12
rect -59 14 -57 18
rect -53 14 -51 18
rect -59 8 -51 14
rect -49 12 -44 18
rect -29 17 -24 33
rect -25 13 -24 17
rect -22 13 -14 33
rect -12 29 -11 33
rect -12 13 -7 29
rect 2 27 7 33
rect 6 23 7 27
rect 9 29 10 33
rect 9 23 14 29
rect -49 8 -48 12
<< pdiffusion >>
rect -62 72 -61 76
rect -66 36 -61 72
rect -59 36 -51 76
rect -49 40 -44 76
rect -25 67 -24 71
rect -29 51 -24 67
rect -22 55 -14 71
rect -22 51 -20 55
rect -16 51 -14 55
rect -12 67 -11 71
rect -12 51 -7 67
rect 6 61 7 65
rect -49 36 -48 40
rect 2 45 7 61
rect 9 49 14 65
rect 9 45 10 49
<< ndcontact >>
rect -66 8 -62 12
rect -57 14 -53 18
rect -29 13 -25 17
rect -11 29 -7 33
rect 2 23 6 27
rect 10 29 14 33
rect -48 8 -44 12
<< pdcontact >>
rect -66 72 -62 76
rect -29 67 -25 71
rect -20 51 -16 55
rect -11 67 -7 71
rect 2 61 6 65
rect -48 36 -44 40
rect 10 45 14 49
<< polysilicon >>
rect -61 76 -59 79
rect -51 76 -49 79
rect -24 71 -22 75
rect -14 71 -12 75
rect 7 65 9 69
rect -61 18 -59 36
rect -51 18 -49 36
rect -24 33 -22 51
rect -14 33 -12 51
rect 7 33 9 45
rect 7 19 9 23
rect -24 9 -22 13
rect -14 9 -12 13
rect -61 5 -59 8
rect -51 5 -49 8
<< polycontact >>
rect -28 40 -24 44
rect -65 19 -61 23
rect -55 25 -51 29
rect -18 34 -14 38
rect 3 34 7 38
<< metal1 >>
rect -72 83 -32 86
rect -66 76 -63 83
rect -35 81 -32 83
rect -35 78 5 81
rect -29 71 -26 78
rect -11 71 -7 78
rect 2 65 5 78
rect -19 50 -16 51
rect -19 47 -7 50
rect -35 41 -28 44
rect -10 38 -7 47
rect 11 38 14 45
rect -72 26 -55 29
rect -47 27 -44 36
rect -35 34 -18 37
rect -10 35 3 38
rect -35 27 -32 34
rect -10 33 -7 35
rect 11 35 18 38
rect 11 33 14 35
rect -47 24 -32 27
rect -72 20 -65 23
rect -47 22 -44 24
rect -56 19 -44 22
rect -56 18 -53 19
rect -29 8 -26 13
rect 2 8 5 23
rect -66 4 -63 8
rect -47 4 -44 8
rect -35 5 5 8
rect -35 4 -32 5
rect -72 1 -32 4
<< labels >>
rlabel metal1 -65 84 -65 85 5 vdd
rlabel metal1 -55 3 -55 3 1 gnd
rlabel metal1 -70 26 -66 28 3 p3_inv
rlabel metal1 -71 21 -69 22 3 p2_inv
rlabel metal1 -41 24 -40 26 7 temp109
rlabel metal1 -23 79 -23 79 5 vdd
rlabel metal1 -14 6 -14 6 1 gnd
rlabel metal1 -33 41 -30 44 1 temp101
rlabel metal1 12 36 14 38 1 p4
<< end >>
