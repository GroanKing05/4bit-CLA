magic
tech scmos
timestamp 1731422623
<< nwell >>
rect 418 -140 450 -121
rect 418 -146 472 -140
rect 420 -174 472 -146
rect 490 -156 567 -134
rect 490 -166 585 -156
rect 122 -195 156 -175
rect 88 -227 156 -195
rect 162 -197 220 -175
rect 162 -207 269 -197
rect 335 -201 369 -181
rect 397 -194 431 -188
rect 186 -227 269 -207
rect 214 -229 269 -227
rect 301 -233 369 -201
rect 375 -220 431 -194
rect 375 -226 400 -220
rect 448 -234 482 -182
rect 533 -186 585 -166
rect 561 -188 585 -186
rect 623 -203 657 -183
rect 688 -188 765 -166
rect 805 -172 837 -153
rect 589 -235 657 -203
rect 670 -198 765 -188
rect 783 -178 837 -172
rect 670 -218 722 -198
rect 783 -206 835 -178
rect 670 -220 694 -218
rect 773 -266 807 -214
rect 824 -226 858 -220
rect 824 -252 880 -226
rect 855 -258 880 -252
rect 30 -314 63 -282
rect 70 -319 102 -293
rect 147 -319 179 -293
rect 186 -314 219 -282
rect 243 -320 276 -288
rect 283 -325 315 -299
rect 360 -325 392 -299
rect 399 -320 432 -288
rect 531 -322 564 -290
rect 571 -327 603 -301
rect 648 -327 680 -301
rect 687 -322 720 -290
<< ntransistor >>
rect 402 -135 412 -133
rect 398 -153 408 -151
rect 398 -163 408 -161
rect 173 -223 175 -213
rect 99 -259 101 -239
rect 109 -259 111 -239
rect 133 -249 135 -239
rect 143 -249 145 -239
rect 197 -249 199 -239
rect 207 -249 209 -239
rect 225 -245 227 -235
rect 246 -261 248 -241
rect 256 -261 258 -241
rect 501 -198 503 -178
rect 511 -198 513 -178
rect 843 -167 853 -165
rect 544 -208 546 -198
rect 554 -208 556 -198
rect 572 -204 574 -194
rect 387 -242 389 -232
rect 312 -265 314 -245
rect 322 -265 324 -245
rect 346 -255 348 -245
rect 356 -255 358 -245
rect 408 -252 410 -232
rect 418 -252 420 -232
rect 847 -185 857 -183
rect 847 -195 857 -193
rect 459 -256 461 -246
rect 469 -256 471 -246
rect 681 -236 683 -226
rect 742 -230 744 -210
rect 752 -230 754 -210
rect 699 -240 701 -230
rect 709 -240 711 -230
rect 600 -267 602 -247
rect 610 -267 612 -247
rect 634 -257 636 -247
rect 644 -257 646 -247
rect 108 -307 118 -305
rect 131 -307 141 -305
rect 321 -313 331 -311
rect 344 -313 354 -311
rect 41 -331 43 -321
rect 50 -331 52 -321
rect 197 -331 199 -321
rect 206 -331 208 -321
rect 784 -288 786 -278
rect 794 -288 796 -278
rect 835 -284 837 -264
rect 845 -284 847 -264
rect 866 -274 868 -264
rect 609 -315 619 -313
rect 632 -315 642 -313
rect 254 -337 256 -327
rect 263 -337 265 -327
rect 410 -337 412 -327
rect 419 -337 421 -327
rect 542 -339 544 -329
rect 551 -339 553 -329
rect 698 -339 700 -329
rect 707 -339 709 -329
<< ptransistor >>
rect 424 -135 444 -133
rect 426 -153 466 -151
rect 501 -160 503 -140
rect 511 -160 513 -140
rect 426 -163 466 -161
rect 99 -221 101 -201
rect 109 -221 111 -201
rect 133 -221 135 -181
rect 143 -221 145 -181
rect 173 -201 175 -181
rect 197 -221 199 -181
rect 207 -221 209 -181
rect 225 -223 227 -203
rect 246 -223 248 -203
rect 256 -223 258 -203
rect 312 -227 314 -207
rect 322 -227 324 -207
rect 346 -227 348 -187
rect 356 -227 358 -187
rect 387 -220 389 -200
rect 408 -214 410 -194
rect 418 -214 420 -194
rect 459 -228 461 -188
rect 469 -228 471 -188
rect 544 -180 546 -140
rect 554 -180 556 -140
rect 572 -182 574 -162
rect 811 -167 831 -165
rect 600 -229 602 -209
rect 610 -229 612 -209
rect 634 -229 636 -189
rect 644 -229 646 -189
rect 681 -214 683 -194
rect 699 -212 701 -172
rect 709 -212 711 -172
rect 742 -192 744 -172
rect 752 -192 754 -172
rect 789 -185 829 -183
rect 789 -195 829 -193
rect 784 -260 786 -220
rect 794 -260 796 -220
rect 835 -246 837 -226
rect 845 -246 847 -226
rect 866 -252 868 -232
rect 41 -308 43 -288
rect 50 -308 52 -288
rect 76 -307 96 -305
rect 153 -307 173 -305
rect 197 -308 199 -288
rect 206 -308 208 -288
rect 254 -314 256 -294
rect 263 -314 265 -294
rect 289 -313 309 -311
rect 366 -313 386 -311
rect 410 -314 412 -294
rect 419 -314 421 -294
rect 542 -316 544 -296
rect 551 -316 553 -296
rect 577 -315 597 -313
rect 654 -315 674 -313
rect 698 -316 700 -296
rect 707 -316 709 -296
<< ndiffusion >>
rect 402 -132 408 -128
rect 402 -133 412 -132
rect 402 -136 412 -135
rect 406 -140 412 -136
rect 402 -150 408 -146
rect 398 -151 408 -150
rect 398 -155 408 -153
rect 398 -159 404 -155
rect 398 -161 408 -159
rect 398 -164 408 -163
rect 402 -168 408 -164
rect 168 -219 173 -213
rect 172 -223 173 -219
rect 175 -217 176 -213
rect 175 -223 180 -217
rect 98 -243 99 -239
rect 94 -259 99 -243
rect 101 -259 109 -239
rect 111 -255 116 -239
rect 128 -245 133 -239
rect 132 -249 133 -245
rect 135 -243 137 -239
rect 141 -243 143 -239
rect 135 -249 143 -243
rect 145 -245 150 -239
rect 145 -249 146 -245
rect 192 -245 197 -239
rect 196 -249 197 -245
rect 199 -243 201 -239
rect 205 -243 207 -239
rect 199 -249 207 -243
rect 209 -245 214 -239
rect 220 -241 225 -235
rect 224 -245 225 -241
rect 227 -239 228 -235
rect 227 -245 232 -239
rect 209 -249 210 -245
rect 111 -259 112 -255
rect 241 -257 246 -241
rect 245 -261 246 -257
rect 248 -261 256 -241
rect 258 -245 259 -241
rect 496 -194 501 -178
rect 500 -198 501 -194
rect 503 -198 511 -178
rect 513 -182 514 -178
rect 513 -198 518 -182
rect 847 -164 853 -160
rect 843 -165 853 -164
rect 843 -168 853 -167
rect 843 -172 849 -168
rect 539 -204 544 -198
rect 543 -208 544 -204
rect 546 -202 548 -198
rect 552 -202 554 -198
rect 546 -208 554 -202
rect 556 -204 561 -198
rect 567 -200 572 -194
rect 571 -204 572 -200
rect 574 -198 575 -194
rect 574 -204 579 -198
rect 556 -208 557 -204
rect 386 -236 387 -232
rect 382 -242 387 -236
rect 389 -238 394 -232
rect 389 -242 390 -238
rect 407 -236 408 -232
rect 258 -261 263 -245
rect 311 -249 312 -245
rect 307 -265 312 -249
rect 314 -265 322 -245
rect 324 -261 329 -245
rect 341 -251 346 -245
rect 345 -255 346 -251
rect 348 -249 350 -245
rect 354 -249 356 -245
rect 348 -255 356 -249
rect 358 -251 363 -245
rect 358 -255 359 -251
rect 403 -252 408 -236
rect 410 -252 418 -232
rect 420 -248 425 -232
rect 847 -182 853 -178
rect 847 -183 857 -182
rect 847 -187 857 -185
rect 851 -191 857 -187
rect 847 -193 857 -191
rect 847 -196 857 -195
rect 847 -200 853 -196
rect 420 -252 421 -248
rect 454 -252 459 -246
rect 458 -256 459 -252
rect 461 -250 463 -246
rect 467 -250 469 -246
rect 461 -256 469 -250
rect 471 -252 476 -246
rect 680 -230 681 -226
rect 676 -236 681 -230
rect 683 -232 688 -226
rect 741 -214 742 -210
rect 737 -230 742 -214
rect 744 -230 752 -210
rect 754 -226 759 -210
rect 754 -230 755 -226
rect 683 -236 684 -232
rect 694 -236 699 -230
rect 698 -240 699 -236
rect 701 -234 703 -230
rect 707 -234 709 -230
rect 701 -240 709 -234
rect 711 -236 716 -230
rect 711 -240 712 -236
rect 471 -256 472 -252
rect 599 -251 600 -247
rect 324 -265 325 -261
rect 595 -267 600 -251
rect 602 -267 610 -247
rect 612 -263 617 -247
rect 629 -253 634 -247
rect 633 -257 634 -253
rect 636 -251 638 -247
rect 642 -251 644 -247
rect 636 -257 644 -251
rect 646 -253 651 -247
rect 646 -257 647 -253
rect 612 -267 613 -263
rect 108 -304 114 -300
rect 108 -305 118 -304
rect 138 -304 141 -300
rect 131 -305 141 -304
rect 108 -308 118 -307
rect 112 -312 118 -308
rect 131 -308 141 -307
rect 131 -312 137 -308
rect 779 -284 784 -278
rect 321 -310 327 -306
rect 321 -311 331 -310
rect 351 -310 354 -306
rect 344 -311 354 -310
rect 40 -325 41 -321
rect 36 -331 41 -325
rect 43 -325 45 -321
rect 49 -325 50 -321
rect 43 -331 50 -325
rect 52 -327 57 -321
rect 52 -331 53 -327
rect 192 -327 197 -321
rect 196 -331 197 -327
rect 199 -325 200 -321
rect 204 -325 206 -321
rect 199 -331 206 -325
rect 208 -325 209 -321
rect 208 -331 213 -325
rect 321 -314 331 -313
rect 325 -318 331 -314
rect 344 -314 354 -313
rect 344 -318 350 -314
rect 783 -288 784 -284
rect 786 -282 788 -278
rect 792 -282 794 -278
rect 786 -288 794 -282
rect 796 -284 801 -278
rect 830 -280 835 -264
rect 834 -284 835 -280
rect 837 -284 845 -264
rect 847 -268 848 -264
rect 847 -284 852 -268
rect 861 -270 866 -264
rect 865 -274 866 -270
rect 868 -268 869 -264
rect 868 -274 873 -268
rect 796 -288 797 -284
rect 609 -312 615 -308
rect 609 -313 619 -312
rect 639 -312 642 -308
rect 632 -313 642 -312
rect 253 -331 254 -327
rect 249 -337 254 -331
rect 256 -331 258 -327
rect 262 -331 263 -327
rect 256 -337 263 -331
rect 265 -333 270 -327
rect 265 -337 266 -333
rect 405 -333 410 -327
rect 409 -337 410 -333
rect 412 -331 413 -327
rect 417 -331 419 -327
rect 412 -337 419 -331
rect 421 -331 422 -327
rect 609 -316 619 -315
rect 613 -320 619 -316
rect 632 -316 642 -315
rect 632 -320 638 -316
rect 421 -337 426 -331
rect 541 -333 542 -329
rect 537 -339 542 -333
rect 544 -333 546 -329
rect 550 -333 551 -329
rect 544 -339 551 -333
rect 553 -335 558 -329
rect 553 -339 554 -335
rect 693 -335 698 -329
rect 697 -339 698 -335
rect 700 -333 701 -329
rect 705 -333 707 -329
rect 700 -339 707 -333
rect 709 -333 710 -329
rect 709 -339 714 -333
<< pdiffusion >>
rect 428 -132 444 -128
rect 424 -133 444 -132
rect 424 -136 444 -135
rect 424 -140 440 -136
rect 500 -144 501 -140
rect 430 -150 466 -146
rect 426 -151 466 -150
rect 426 -161 466 -153
rect 496 -160 501 -144
rect 503 -156 511 -140
rect 503 -160 505 -156
rect 509 -160 511 -156
rect 513 -144 514 -140
rect 513 -160 518 -144
rect 543 -144 544 -140
rect 426 -164 466 -163
rect 426 -168 462 -164
rect 132 -185 133 -181
rect 98 -205 99 -201
rect 94 -221 99 -205
rect 101 -217 109 -201
rect 101 -221 103 -217
rect 107 -221 109 -217
rect 111 -205 112 -201
rect 111 -221 116 -205
rect 128 -221 133 -185
rect 135 -221 143 -181
rect 145 -217 150 -181
rect 172 -185 173 -181
rect 168 -201 173 -185
rect 175 -197 180 -181
rect 175 -201 176 -197
rect 196 -185 197 -181
rect 145 -221 146 -217
rect 192 -221 197 -185
rect 199 -221 207 -181
rect 209 -217 214 -181
rect 345 -191 346 -187
rect 209 -221 210 -217
rect 224 -207 225 -203
rect 220 -223 225 -207
rect 227 -219 232 -203
rect 227 -223 228 -219
rect 245 -207 246 -203
rect 241 -223 246 -207
rect 248 -219 256 -203
rect 248 -223 250 -219
rect 254 -223 256 -219
rect 258 -207 259 -203
rect 258 -223 263 -207
rect 311 -211 312 -207
rect 307 -227 312 -211
rect 314 -223 322 -207
rect 314 -227 316 -223
rect 320 -227 322 -223
rect 324 -211 325 -207
rect 324 -227 329 -211
rect 341 -227 346 -191
rect 348 -227 356 -187
rect 358 -223 363 -187
rect 407 -198 408 -194
rect 382 -216 387 -200
rect 386 -220 387 -216
rect 389 -204 390 -200
rect 389 -220 394 -204
rect 403 -214 408 -198
rect 410 -210 418 -194
rect 410 -214 412 -210
rect 416 -214 418 -210
rect 420 -198 421 -194
rect 420 -214 425 -198
rect 358 -227 359 -223
rect 454 -224 459 -188
rect 458 -228 459 -224
rect 461 -228 469 -188
rect 471 -192 472 -188
rect 471 -228 476 -192
rect 539 -180 544 -144
rect 546 -180 554 -140
rect 556 -176 561 -140
rect 556 -180 557 -176
rect 571 -166 572 -162
rect 567 -182 572 -166
rect 574 -178 579 -162
rect 811 -164 827 -160
rect 811 -165 831 -164
rect 811 -168 831 -167
rect 815 -172 831 -168
rect 574 -182 575 -178
rect 633 -193 634 -189
rect 599 -213 600 -209
rect 595 -229 600 -213
rect 602 -225 610 -209
rect 602 -229 604 -225
rect 608 -229 610 -225
rect 612 -213 613 -209
rect 612 -229 617 -213
rect 629 -229 634 -193
rect 636 -229 644 -189
rect 646 -225 651 -189
rect 676 -210 681 -194
rect 680 -214 681 -210
rect 683 -198 684 -194
rect 683 -214 688 -198
rect 694 -208 699 -172
rect 698 -212 699 -208
rect 701 -212 709 -172
rect 711 -176 712 -172
rect 711 -212 716 -176
rect 741 -176 742 -172
rect 737 -192 742 -176
rect 744 -188 752 -172
rect 744 -192 746 -188
rect 750 -192 752 -188
rect 754 -176 755 -172
rect 754 -192 759 -176
rect 789 -182 825 -178
rect 789 -183 829 -182
rect 789 -193 829 -185
rect 789 -196 829 -195
rect 793 -200 829 -196
rect 646 -229 647 -225
rect 783 -224 784 -220
rect 779 -260 784 -224
rect 786 -260 794 -220
rect 796 -256 801 -220
rect 834 -230 835 -226
rect 830 -246 835 -230
rect 837 -242 845 -226
rect 837 -246 839 -242
rect 843 -246 845 -242
rect 847 -230 848 -226
rect 847 -246 852 -230
rect 865 -236 866 -232
rect 796 -260 797 -256
rect 861 -252 866 -236
rect 868 -248 873 -232
rect 868 -252 869 -248
rect 36 -304 41 -288
rect 40 -308 41 -304
rect 43 -302 50 -288
rect 43 -306 45 -302
rect 49 -306 50 -302
rect 43 -308 50 -306
rect 52 -292 53 -288
rect 52 -308 57 -292
rect 196 -292 197 -288
rect 81 -304 96 -299
rect 76 -305 96 -304
rect 153 -304 168 -299
rect 153 -305 173 -304
rect 76 -308 96 -307
rect 76 -312 92 -308
rect 153 -308 173 -307
rect 192 -308 197 -292
rect 199 -302 206 -288
rect 199 -306 200 -302
rect 204 -306 206 -302
rect 199 -308 206 -306
rect 208 -304 213 -288
rect 208 -308 209 -304
rect 157 -312 173 -308
rect 249 -310 254 -294
rect 253 -314 254 -310
rect 256 -308 263 -294
rect 256 -312 258 -308
rect 262 -312 263 -308
rect 256 -314 263 -312
rect 265 -298 266 -294
rect 265 -314 270 -298
rect 409 -298 410 -294
rect 294 -310 309 -305
rect 289 -311 309 -310
rect 366 -310 381 -305
rect 366 -311 386 -310
rect 289 -314 309 -313
rect 289 -318 305 -314
rect 366 -314 386 -313
rect 405 -314 410 -298
rect 412 -308 419 -294
rect 412 -312 413 -308
rect 417 -312 419 -308
rect 412 -314 419 -312
rect 421 -310 426 -294
rect 421 -314 422 -310
rect 537 -312 542 -296
rect 370 -318 386 -314
rect 541 -316 542 -312
rect 544 -310 551 -296
rect 544 -314 546 -310
rect 550 -314 551 -310
rect 544 -316 551 -314
rect 553 -300 554 -296
rect 553 -316 558 -300
rect 697 -300 698 -296
rect 582 -312 597 -307
rect 577 -313 597 -312
rect 654 -312 669 -307
rect 654 -313 674 -312
rect 577 -316 597 -315
rect 577 -320 593 -316
rect 654 -316 674 -315
rect 693 -316 698 -300
rect 700 -310 707 -296
rect 700 -314 701 -310
rect 705 -314 707 -310
rect 700 -316 707 -314
rect 709 -312 714 -296
rect 709 -316 710 -312
rect 658 -320 674 -316
<< ndcontact >>
rect 408 -132 412 -128
rect 402 -140 406 -136
rect 398 -150 402 -146
rect 404 -159 408 -155
rect 398 -168 402 -164
rect 168 -223 172 -219
rect 176 -217 180 -213
rect 94 -243 98 -239
rect 128 -249 132 -245
rect 137 -243 141 -239
rect 146 -249 150 -245
rect 192 -249 196 -245
rect 201 -243 205 -239
rect 220 -245 224 -241
rect 228 -239 232 -235
rect 210 -249 214 -245
rect 112 -259 116 -255
rect 241 -261 245 -257
rect 259 -245 263 -241
rect 496 -198 500 -194
rect 514 -182 518 -178
rect 843 -164 847 -160
rect 849 -172 853 -168
rect 539 -208 543 -204
rect 548 -202 552 -198
rect 567 -204 571 -200
rect 575 -198 579 -194
rect 557 -208 561 -204
rect 382 -236 386 -232
rect 390 -242 394 -238
rect 403 -236 407 -232
rect 307 -249 311 -245
rect 341 -255 345 -251
rect 350 -249 354 -245
rect 359 -255 363 -251
rect 853 -182 857 -178
rect 847 -191 851 -187
rect 853 -200 857 -196
rect 421 -252 425 -248
rect 454 -256 458 -252
rect 463 -250 467 -246
rect 676 -230 680 -226
rect 737 -214 741 -210
rect 755 -230 759 -226
rect 684 -236 688 -232
rect 694 -240 698 -236
rect 703 -234 707 -230
rect 712 -240 716 -236
rect 472 -256 476 -252
rect 595 -251 599 -247
rect 325 -265 329 -261
rect 629 -257 633 -253
rect 638 -251 642 -247
rect 647 -257 651 -253
rect 613 -267 617 -263
rect 114 -304 118 -300
rect 131 -304 138 -300
rect 108 -312 112 -308
rect 137 -312 141 -308
rect 327 -310 331 -306
rect 344 -310 351 -306
rect 36 -325 40 -321
rect 45 -325 49 -321
rect 53 -331 57 -327
rect 192 -331 196 -327
rect 200 -325 204 -321
rect 209 -325 213 -321
rect 321 -318 325 -314
rect 350 -318 354 -314
rect 779 -288 783 -284
rect 788 -282 792 -278
rect 830 -284 834 -280
rect 848 -268 852 -264
rect 861 -274 865 -270
rect 869 -268 873 -264
rect 797 -288 801 -284
rect 615 -312 619 -308
rect 632 -312 639 -308
rect 249 -331 253 -327
rect 258 -331 262 -327
rect 266 -337 270 -333
rect 405 -337 409 -333
rect 413 -331 417 -327
rect 422 -331 426 -327
rect 609 -320 613 -316
rect 638 -320 642 -316
rect 537 -333 541 -329
rect 546 -333 550 -329
rect 554 -339 558 -335
rect 693 -339 697 -335
rect 701 -333 705 -329
rect 710 -333 714 -329
<< pdcontact >>
rect 424 -132 428 -128
rect 440 -140 444 -136
rect 496 -144 500 -140
rect 426 -150 430 -146
rect 505 -160 509 -156
rect 514 -144 518 -140
rect 539 -144 543 -140
rect 462 -168 466 -164
rect 128 -185 132 -181
rect 94 -205 98 -201
rect 103 -221 107 -217
rect 112 -205 116 -201
rect 168 -185 172 -181
rect 176 -201 180 -197
rect 192 -185 196 -181
rect 146 -221 150 -217
rect 341 -191 345 -187
rect 210 -221 214 -217
rect 220 -207 224 -203
rect 228 -223 232 -219
rect 241 -207 245 -203
rect 250 -223 254 -219
rect 259 -207 263 -203
rect 307 -211 311 -207
rect 316 -227 320 -223
rect 325 -211 329 -207
rect 403 -198 407 -194
rect 382 -220 386 -216
rect 390 -204 394 -200
rect 412 -214 416 -210
rect 421 -198 425 -194
rect 359 -227 363 -223
rect 454 -228 458 -224
rect 472 -192 476 -188
rect 557 -180 561 -176
rect 567 -166 571 -162
rect 827 -164 831 -160
rect 811 -172 815 -168
rect 575 -182 579 -178
rect 629 -193 633 -189
rect 595 -213 599 -209
rect 604 -229 608 -225
rect 613 -213 617 -209
rect 676 -214 680 -210
rect 684 -198 688 -194
rect 694 -212 698 -208
rect 712 -176 716 -172
rect 737 -176 741 -172
rect 746 -192 750 -188
rect 755 -176 759 -172
rect 825 -182 829 -178
rect 789 -200 793 -196
rect 647 -229 651 -225
rect 779 -224 783 -220
rect 830 -230 834 -226
rect 839 -246 843 -242
rect 848 -230 852 -226
rect 861 -236 865 -232
rect 797 -260 801 -256
rect 869 -252 873 -248
rect 36 -308 40 -304
rect 45 -306 49 -302
rect 53 -292 57 -288
rect 192 -292 196 -288
rect 92 -312 96 -308
rect 200 -306 204 -302
rect 209 -308 213 -304
rect 153 -312 157 -308
rect 249 -314 253 -310
rect 258 -312 262 -308
rect 266 -298 270 -294
rect 405 -298 409 -294
rect 305 -318 309 -314
rect 413 -312 417 -308
rect 422 -314 426 -310
rect 366 -318 370 -314
rect 537 -316 541 -312
rect 546 -314 550 -310
rect 554 -300 558 -296
rect 693 -300 697 -296
rect 593 -320 597 -316
rect 701 -314 705 -310
rect 710 -316 714 -312
rect 654 -320 658 -316
<< polysilicon >>
rect 399 -135 402 -133
rect 412 -135 424 -133
rect 444 -135 447 -133
rect 501 -140 503 -136
rect 511 -140 513 -136
rect 544 -140 546 -137
rect 554 -140 556 -137
rect 395 -153 398 -151
rect 408 -153 426 -151
rect 466 -153 469 -151
rect 395 -163 398 -161
rect 408 -163 426 -161
rect 466 -163 469 -161
rect 133 -181 135 -178
rect 143 -181 145 -178
rect 173 -181 175 -177
rect 501 -178 503 -160
rect 511 -178 513 -160
rect 197 -181 199 -178
rect 207 -181 209 -178
rect 99 -201 101 -197
rect 109 -201 111 -197
rect 173 -213 175 -201
rect 99 -239 101 -221
rect 109 -239 111 -221
rect 133 -239 135 -221
rect 143 -239 145 -221
rect 346 -187 348 -184
rect 356 -187 358 -184
rect 225 -203 227 -200
rect 246 -203 248 -199
rect 256 -203 258 -199
rect 173 -227 175 -223
rect 197 -239 199 -221
rect 207 -239 209 -221
rect 312 -207 314 -203
rect 322 -207 324 -203
rect 225 -235 227 -223
rect 246 -241 248 -223
rect 256 -241 258 -223
rect 459 -188 461 -185
rect 469 -188 471 -185
rect 408 -194 410 -190
rect 418 -194 420 -190
rect 387 -200 389 -196
rect 225 -248 227 -245
rect 133 -252 135 -249
rect 143 -252 145 -249
rect 197 -252 199 -249
rect 207 -252 209 -249
rect 99 -263 101 -259
rect 109 -263 111 -259
rect 312 -245 314 -227
rect 322 -245 324 -227
rect 346 -245 348 -227
rect 356 -245 358 -227
rect 387 -232 389 -220
rect 408 -232 410 -214
rect 418 -232 420 -214
rect 572 -162 574 -159
rect 544 -198 546 -180
rect 554 -198 556 -180
rect 808 -167 811 -165
rect 831 -167 843 -165
rect 853 -167 856 -165
rect 699 -172 701 -169
rect 709 -172 711 -169
rect 742 -172 744 -168
rect 752 -172 754 -168
rect 572 -194 574 -182
rect 634 -189 636 -186
rect 644 -189 646 -186
rect 501 -202 503 -198
rect 511 -202 513 -198
rect 572 -207 574 -204
rect 544 -211 546 -208
rect 554 -211 556 -208
rect 600 -209 602 -205
rect 610 -209 612 -205
rect 246 -265 248 -261
rect 256 -265 258 -261
rect 387 -246 389 -242
rect 459 -246 461 -228
rect 469 -246 471 -228
rect 681 -194 683 -191
rect 786 -185 789 -183
rect 829 -185 847 -183
rect 857 -185 860 -183
rect 742 -210 744 -192
rect 752 -210 754 -192
rect 786 -195 789 -193
rect 829 -195 847 -193
rect 857 -195 860 -193
rect 681 -226 683 -214
rect 346 -258 348 -255
rect 356 -258 358 -255
rect 408 -256 410 -252
rect 418 -256 420 -252
rect 600 -247 602 -229
rect 610 -247 612 -229
rect 634 -247 636 -229
rect 644 -247 646 -229
rect 699 -230 701 -212
rect 709 -230 711 -212
rect 784 -220 786 -217
rect 794 -220 796 -217
rect 681 -239 683 -236
rect 742 -234 744 -230
rect 752 -234 754 -230
rect 699 -243 701 -240
rect 709 -243 711 -240
rect 459 -259 461 -256
rect 469 -259 471 -256
rect 312 -269 314 -265
rect 322 -269 324 -265
rect 634 -260 636 -257
rect 644 -260 646 -257
rect 835 -226 837 -222
rect 845 -226 847 -222
rect 866 -232 868 -228
rect 600 -271 602 -267
rect 610 -271 612 -267
rect 41 -288 43 -276
rect 50 -288 52 -285
rect 197 -288 199 -285
rect 206 -288 208 -276
rect 784 -278 786 -260
rect 794 -278 796 -260
rect 835 -264 837 -246
rect 845 -264 847 -246
rect 866 -264 868 -252
rect 72 -307 76 -305
rect 96 -307 108 -305
rect 118 -307 122 -305
rect 127 -307 131 -305
rect 141 -307 153 -305
rect 173 -307 177 -305
rect 41 -314 43 -308
rect 41 -321 43 -317
rect 50 -321 52 -308
rect 254 -294 256 -282
rect 263 -294 265 -291
rect 410 -294 412 -291
rect 419 -294 421 -282
rect 197 -321 199 -308
rect 206 -314 208 -308
rect 285 -313 289 -311
rect 309 -313 321 -311
rect 331 -313 335 -311
rect 340 -313 344 -311
rect 354 -313 366 -311
rect 386 -313 390 -311
rect 206 -321 208 -317
rect 254 -320 256 -314
rect 254 -327 256 -323
rect 263 -327 265 -314
rect 542 -296 544 -284
rect 551 -296 553 -293
rect 698 -296 700 -293
rect 707 -296 709 -284
rect 866 -278 868 -274
rect 835 -288 837 -284
rect 845 -288 847 -284
rect 784 -291 786 -288
rect 794 -291 796 -288
rect 410 -327 412 -314
rect 419 -320 421 -314
rect 573 -315 577 -313
rect 597 -315 609 -313
rect 619 -315 623 -313
rect 628 -315 632 -313
rect 642 -315 654 -313
rect 674 -315 678 -313
rect 542 -322 544 -316
rect 419 -327 421 -323
rect 41 -333 43 -331
rect 41 -337 42 -333
rect 50 -334 52 -331
rect 197 -334 199 -331
rect 206 -333 208 -331
rect 207 -337 208 -333
rect 542 -329 544 -325
rect 551 -329 553 -316
rect 698 -329 700 -316
rect 707 -322 709 -316
rect 707 -329 709 -325
rect 41 -338 43 -337
rect 206 -338 208 -337
rect 254 -339 256 -337
rect 254 -343 255 -339
rect 263 -340 265 -337
rect 410 -340 412 -337
rect 419 -339 421 -337
rect 420 -343 421 -339
rect 254 -344 256 -343
rect 419 -344 421 -343
rect 542 -341 544 -339
rect 542 -345 543 -341
rect 551 -342 553 -339
rect 698 -342 700 -339
rect 707 -341 709 -339
rect 708 -345 709 -341
rect 542 -346 544 -345
rect 707 -346 709 -345
<< polycontact >>
rect 413 -139 417 -135
rect 415 -157 419 -153
rect 409 -167 413 -163
rect 497 -171 501 -167
rect 507 -177 511 -173
rect 169 -212 173 -208
rect 101 -238 105 -234
rect 111 -232 115 -228
rect 129 -238 133 -234
rect 139 -232 143 -228
rect 193 -238 197 -234
rect 203 -232 207 -228
rect 221 -234 225 -230
rect 242 -234 246 -230
rect 252 -240 256 -236
rect 314 -244 318 -240
rect 324 -238 328 -234
rect 342 -244 346 -240
rect 352 -238 356 -234
rect 389 -231 393 -227
rect 410 -231 414 -227
rect 420 -225 424 -221
rect 540 -197 544 -193
rect 550 -191 554 -187
rect 838 -171 842 -167
rect 568 -193 572 -189
rect 461 -239 465 -235
rect 744 -209 748 -205
rect 836 -189 840 -185
rect 754 -203 758 -199
rect 842 -199 846 -195
rect 683 -225 687 -221
rect 471 -245 475 -241
rect 602 -246 606 -242
rect 612 -240 616 -236
rect 630 -246 634 -242
rect 640 -240 644 -236
rect 701 -223 705 -219
rect 711 -229 715 -225
rect 831 -257 835 -253
rect 43 -281 47 -277
rect 202 -281 206 -277
rect 780 -277 784 -273
rect 790 -271 794 -267
rect 841 -263 845 -259
rect 862 -263 866 -259
rect 103 -305 107 -301
rect 142 -305 146 -301
rect 256 -287 260 -283
rect 415 -287 419 -283
rect 52 -319 56 -315
rect 193 -319 197 -315
rect 316 -311 320 -307
rect 355 -311 359 -307
rect 544 -289 548 -285
rect 703 -289 707 -285
rect 265 -325 269 -321
rect 406 -325 410 -321
rect 604 -313 608 -309
rect 643 -313 647 -309
rect 42 -337 46 -333
rect 203 -337 207 -333
rect 553 -327 557 -323
rect 694 -327 698 -323
rect 255 -343 259 -339
rect 416 -343 420 -339
rect 543 -345 547 -341
rect 704 -345 708 -341
<< metal1 >>
rect 414 -124 454 -121
rect 414 -128 417 -124
rect 412 -131 424 -128
rect 451 -130 454 -124
rect 451 -133 482 -130
rect 495 -133 570 -130
rect 391 -140 402 -137
rect 391 -146 394 -140
rect 414 -146 417 -139
rect 444 -140 471 -137
rect 391 -149 398 -146
rect 391 -164 394 -149
rect 409 -149 426 -146
rect 409 -155 412 -149
rect 408 -158 412 -155
rect 119 -172 122 -171
rect 394 -168 398 -165
rect 127 -172 223 -171
rect 409 -172 413 -167
rect 119 -174 223 -172
rect 119 -191 122 -174
rect 128 -181 131 -174
rect 168 -181 171 -174
rect 192 -181 195 -174
rect 88 -194 122 -191
rect 220 -193 223 -174
rect 332 -178 335 -177
rect 416 -174 419 -157
rect 473 -165 476 -142
rect 466 -168 476 -165
rect 340 -178 397 -177
rect 332 -180 397 -178
rect 473 -178 476 -168
rect 479 -167 482 -133
rect 496 -140 499 -133
rect 514 -140 518 -133
rect 539 -140 542 -133
rect 567 -152 570 -133
rect 567 -155 590 -152
rect 506 -161 509 -160
rect 506 -164 518 -161
rect 479 -170 497 -167
rect 515 -173 518 -164
rect 567 -162 570 -155
rect 494 -177 507 -174
rect 515 -176 536 -173
rect 587 -174 590 -155
rect 801 -156 841 -153
rect 685 -165 760 -162
rect 801 -162 804 -156
rect 838 -160 841 -156
rect 773 -165 804 -162
rect 831 -163 843 -160
rect 587 -175 628 -174
rect 515 -178 518 -176
rect 94 -201 98 -194
rect 113 -201 116 -194
rect 220 -196 269 -193
rect 177 -208 180 -201
rect 220 -203 223 -196
rect 241 -203 244 -196
rect 259 -203 263 -196
rect 332 -197 335 -180
rect 341 -187 344 -180
rect 394 -184 397 -180
rect 428 -181 476 -178
rect 428 -184 431 -181
rect 391 -187 431 -184
rect 301 -200 335 -197
rect 391 -200 394 -187
rect 403 -194 407 -187
rect 422 -194 425 -187
rect 473 -188 476 -181
rect 533 -187 536 -176
rect 587 -177 623 -175
rect 533 -190 550 -187
rect 558 -189 561 -180
rect 576 -189 579 -182
rect 620 -180 623 -177
rect 628 -180 657 -179
rect 620 -182 657 -180
rect 558 -192 568 -189
rect 536 -196 540 -193
rect 558 -194 561 -192
rect 576 -192 586 -189
rect 576 -194 579 -192
rect 549 -197 561 -194
rect 549 -198 552 -197
rect 307 -207 311 -200
rect 326 -207 329 -200
rect 496 -203 499 -198
rect 620 -199 623 -182
rect 629 -189 632 -182
rect 685 -194 688 -165
rect 713 -172 716 -165
rect 737 -172 741 -165
rect 756 -172 759 -165
rect 746 -193 749 -192
rect 737 -196 749 -193
rect 162 -211 169 -208
rect 103 -222 106 -221
rect 94 -225 106 -222
rect 94 -234 97 -225
rect 115 -231 139 -228
rect 147 -230 150 -221
rect 147 -233 153 -230
rect 75 -237 97 -234
rect 94 -239 97 -237
rect 105 -238 129 -235
rect 147 -235 150 -233
rect 138 -238 150 -235
rect 162 -235 165 -211
rect 177 -211 188 -208
rect 487 -206 535 -203
rect 589 -202 623 -199
rect 177 -213 180 -211
rect 168 -228 171 -223
rect 185 -228 188 -211
rect 412 -215 415 -214
rect 168 -231 181 -228
rect 185 -231 203 -228
rect 162 -238 174 -235
rect 120 -239 125 -238
rect 138 -239 141 -238
rect 87 -263 90 -246
rect 128 -253 131 -249
rect 147 -252 150 -249
rect 75 -266 90 -263
rect 113 -264 116 -259
rect 119 -256 147 -253
rect 119 -264 122 -256
rect 75 -278 78 -266
rect 113 -267 122 -264
rect 47 -281 78 -278
rect 66 -288 69 -281
rect 57 -291 106 -288
rect 123 -291 126 -275
rect 37 -315 40 -308
rect 103 -301 106 -291
rect 121 -295 128 -291
rect 136 -300 139 -256
rect 171 -259 174 -238
rect 178 -251 181 -231
rect 211 -230 214 -221
rect 403 -218 415 -215
rect 229 -230 232 -223
rect 251 -224 254 -223
rect 251 -227 263 -224
rect 211 -233 221 -230
rect 190 -237 193 -234
rect 211 -235 214 -233
rect 229 -233 242 -230
rect 229 -235 232 -233
rect 202 -238 214 -235
rect 202 -239 205 -238
rect 260 -236 263 -227
rect 382 -227 385 -220
rect 403 -227 406 -218
rect 424 -224 451 -221
rect 316 -228 319 -227
rect 307 -231 319 -228
rect 240 -240 252 -237
rect 260 -239 269 -236
rect 260 -241 263 -239
rect 192 -253 195 -249
rect 211 -253 214 -249
rect 220 -252 223 -245
rect 182 -256 219 -253
rect 266 -257 269 -239
rect 171 -262 186 -259
rect 183 -268 186 -262
rect 266 -260 282 -257
rect 241 -265 244 -261
rect 293 -263 296 -233
rect 307 -240 310 -231
rect 328 -237 352 -234
rect 360 -236 363 -227
rect 379 -230 385 -227
rect 382 -232 385 -230
rect 393 -230 406 -227
rect 403 -232 406 -230
rect 414 -231 433 -228
rect 360 -239 372 -236
rect 448 -237 451 -224
rect 454 -237 457 -228
rect 304 -243 310 -240
rect 307 -245 310 -243
rect 318 -244 342 -241
rect 360 -241 363 -239
rect 351 -244 363 -241
rect 369 -242 372 -239
rect 448 -240 457 -237
rect 465 -238 478 -235
rect 333 -245 338 -244
rect 351 -245 354 -244
rect 276 -266 296 -263
rect 245 -269 266 -266
rect 276 -274 279 -266
rect 300 -269 303 -252
rect 341 -259 344 -255
rect 360 -257 363 -255
rect 391 -256 394 -242
rect 454 -242 457 -240
rect 454 -245 466 -242
rect 475 -244 483 -241
rect 463 -246 466 -245
rect 360 -259 390 -257
rect 332 -260 390 -259
rect 288 -272 303 -269
rect 326 -270 329 -265
rect 332 -262 363 -260
rect 422 -257 425 -252
rect 395 -260 431 -257
rect 454 -260 457 -256
rect 473 -260 476 -256
rect 487 -260 490 -206
rect 532 -212 535 -206
rect 539 -212 542 -208
rect 558 -212 561 -208
rect 567 -212 570 -204
rect 532 -215 570 -212
rect 595 -209 599 -202
rect 614 -209 617 -202
rect 737 -205 740 -196
rect 773 -199 776 -165
rect 758 -202 776 -199
rect 784 -172 811 -169
rect 779 -197 782 -174
rect 838 -178 841 -171
rect 853 -172 864 -169
rect 861 -178 864 -172
rect 829 -181 846 -178
rect 843 -187 846 -181
rect 857 -181 864 -178
rect 779 -200 789 -197
rect 719 -208 740 -205
rect 332 -270 335 -262
rect 169 -280 170 -275
rect 175 -278 176 -275
rect 175 -280 202 -278
rect 169 -281 202 -280
rect 169 -282 176 -281
rect 180 -288 183 -281
rect 288 -284 291 -272
rect 326 -273 335 -270
rect 260 -287 291 -284
rect 118 -303 131 -300
rect 138 -304 139 -300
rect 143 -291 192 -288
rect 143 -301 146 -291
rect 279 -294 282 -287
rect 270 -297 319 -294
rect 336 -297 339 -281
rect 45 -309 48 -306
rect 96 -312 108 -309
rect 141 -312 153 -309
rect 201 -309 204 -306
rect 28 -317 40 -315
rect 33 -318 40 -317
rect 37 -321 40 -318
rect 45 -321 48 -314
rect 56 -319 62 -316
rect 103 -320 106 -312
rect 73 -323 106 -320
rect 143 -320 146 -312
rect 187 -319 193 -316
rect 143 -323 176 -320
rect 201 -321 204 -314
rect 73 -326 76 -323
rect 60 -328 76 -326
rect 57 -329 76 -328
rect 173 -326 176 -323
rect 209 -315 212 -308
rect 209 -317 221 -315
rect 209 -318 216 -317
rect 209 -321 212 -318
rect 250 -321 253 -314
rect 316 -307 319 -297
rect 334 -301 341 -297
rect 349 -306 352 -262
rect 427 -263 490 -260
rect 567 -257 570 -215
rect 676 -221 679 -214
rect 694 -221 697 -212
rect 719 -219 722 -208
rect 737 -210 740 -208
rect 748 -209 762 -206
rect 779 -210 782 -200
rect 836 -206 839 -189
rect 843 -190 847 -187
rect 861 -196 864 -181
rect 842 -202 846 -199
rect 857 -200 861 -197
rect 779 -213 827 -210
rect 669 -224 679 -221
rect 604 -230 607 -229
rect 595 -233 607 -230
rect 581 -265 584 -235
rect 595 -240 598 -233
rect 616 -239 640 -236
rect 648 -238 651 -229
rect 676 -226 679 -224
rect 687 -224 697 -221
rect 705 -222 722 -219
rect 779 -220 782 -213
rect 824 -216 827 -213
rect 824 -219 864 -216
rect 694 -226 697 -224
rect 694 -229 706 -226
rect 715 -228 719 -225
rect 703 -230 706 -229
rect 830 -226 833 -219
rect 848 -226 852 -219
rect 756 -235 759 -230
rect 861 -232 864 -219
rect 594 -245 598 -240
rect 648 -241 660 -238
rect 595 -247 598 -245
rect 606 -246 630 -243
rect 648 -243 651 -241
rect 639 -246 651 -243
rect 657 -243 660 -241
rect 621 -247 626 -246
rect 639 -247 642 -246
rect 685 -244 688 -236
rect 694 -244 697 -240
rect 713 -244 716 -240
rect 720 -238 768 -235
rect 720 -244 723 -238
rect 685 -247 723 -244
rect 564 -268 584 -265
rect 396 -274 399 -272
rect 564 -276 567 -268
rect 588 -271 591 -254
rect 629 -261 632 -257
rect 648 -259 651 -257
rect 648 -261 649 -259
rect 576 -274 591 -271
rect 614 -272 617 -267
rect 620 -264 649 -261
rect 620 -272 623 -264
rect 382 -286 383 -281
rect 388 -284 389 -281
rect 388 -286 415 -284
rect 382 -287 415 -286
rect 382 -288 389 -287
rect 393 -294 396 -287
rect 576 -286 579 -274
rect 614 -275 623 -272
rect 548 -289 579 -286
rect 331 -309 344 -306
rect 351 -310 352 -306
rect 356 -297 405 -294
rect 356 -307 359 -297
rect 567 -296 570 -289
rect 558 -299 607 -296
rect 624 -299 627 -283
rect 258 -315 261 -312
rect 309 -318 321 -315
rect 354 -318 366 -315
rect 414 -315 417 -312
rect 241 -323 253 -321
rect 173 -328 189 -326
rect 173 -329 192 -328
rect 57 -331 63 -329
rect 60 -334 63 -331
rect 46 -337 63 -334
rect 186 -331 192 -329
rect 246 -324 253 -323
rect 250 -327 253 -324
rect 258 -327 261 -320
rect 269 -325 275 -322
rect 316 -326 319 -318
rect 286 -329 319 -326
rect 356 -326 359 -318
rect 400 -325 406 -322
rect 356 -329 389 -326
rect 414 -327 417 -320
rect 186 -334 189 -331
rect 286 -332 289 -329
rect 186 -337 203 -334
rect 273 -334 289 -332
rect 270 -335 289 -334
rect 386 -332 389 -329
rect 422 -321 425 -314
rect 422 -323 434 -321
rect 538 -323 541 -316
rect 604 -309 607 -299
rect 622 -303 629 -299
rect 637 -308 640 -264
rect 670 -288 671 -283
rect 676 -286 677 -283
rect 676 -288 703 -286
rect 670 -289 703 -288
rect 670 -290 677 -289
rect 681 -296 684 -289
rect 765 -292 768 -238
rect 840 -247 843 -246
rect 840 -250 852 -247
rect 804 -256 831 -253
rect 777 -270 790 -267
rect 798 -269 801 -260
rect 804 -269 807 -256
rect 849 -259 852 -250
rect 870 -259 873 -252
rect 828 -263 841 -260
rect 849 -262 862 -259
rect 849 -264 852 -262
rect 870 -262 876 -259
rect 870 -264 873 -262
rect 798 -272 807 -269
rect 772 -276 780 -273
rect 798 -274 801 -272
rect 789 -277 801 -274
rect 789 -278 792 -277
rect 779 -292 782 -288
rect 798 -292 801 -288
rect 830 -289 833 -284
rect 861 -288 864 -274
rect 824 -292 860 -289
rect 765 -295 828 -292
rect 619 -311 632 -308
rect 639 -312 640 -308
rect 644 -299 693 -296
rect 644 -309 647 -299
rect 546 -317 549 -314
rect 597 -320 609 -317
rect 642 -320 654 -317
rect 702 -317 705 -314
rect 422 -324 429 -323
rect 422 -327 425 -324
rect 529 -325 541 -323
rect 534 -326 541 -325
rect 538 -329 541 -326
rect 386 -334 402 -332
rect 546 -329 549 -322
rect 557 -327 563 -324
rect 604 -328 607 -320
rect 574 -331 607 -328
rect 644 -328 647 -320
rect 688 -327 694 -324
rect 644 -331 677 -328
rect 702 -329 705 -322
rect 386 -335 405 -334
rect 270 -337 276 -335
rect 273 -340 276 -337
rect 259 -343 276 -340
rect 399 -337 405 -335
rect 574 -334 577 -331
rect 399 -340 402 -337
rect 561 -336 577 -334
rect 558 -337 577 -336
rect 674 -334 677 -331
rect 710 -323 713 -316
rect 710 -325 722 -323
rect 710 -326 717 -325
rect 710 -329 713 -326
rect 674 -336 690 -334
rect 674 -337 693 -336
rect 558 -339 564 -337
rect 399 -343 416 -340
rect 561 -342 564 -339
rect 547 -345 564 -342
rect 687 -339 693 -337
rect 687 -342 690 -339
rect 687 -345 704 -342
<< m2contact >>
rect 490 -133 495 -128
rect 471 -142 476 -137
rect 407 -177 412 -172
rect 416 -179 421 -174
rect 760 -165 765 -160
rect 79 -227 85 -222
rect 70 -238 75 -233
rect 120 -228 125 -223
rect 153 -234 158 -229
rect 86 -246 91 -241
rect 120 -244 125 -239
rect 62 -273 67 -268
rect 116 -296 121 -291
rect 128 -296 133 -291
rect 147 -257 152 -252
rect 185 -239 190 -234
rect 293 -233 298 -228
rect 235 -242 240 -237
rect 177 -256 182 -251
rect 219 -257 224 -252
rect 282 -260 287 -255
rect 299 -243 304 -238
rect 333 -234 338 -229
rect 374 -232 379 -227
rect 478 -238 483 -233
rect 299 -252 304 -247
rect 333 -250 338 -245
rect 369 -247 374 -242
rect 182 -273 187 -268
rect 240 -270 245 -265
rect 479 -249 484 -244
rect 779 -174 784 -169
rect 275 -279 280 -274
rect 44 -314 49 -309
rect 200 -314 205 -309
rect 329 -302 334 -297
rect 341 -302 346 -297
rect 762 -210 767 -205
rect 834 -211 839 -206
rect 581 -235 586 -230
rect 567 -262 572 -257
rect 621 -236 626 -231
rect 588 -245 594 -240
rect 587 -254 592 -249
rect 621 -252 626 -247
rect 657 -248 662 -243
rect 395 -279 400 -274
rect 649 -264 654 -259
rect 563 -281 568 -276
rect 257 -320 262 -315
rect 413 -320 418 -315
rect 617 -304 622 -299
rect 629 -304 634 -299
rect 683 -281 688 -276
rect 772 -270 777 -265
rect 876 -264 881 -259
rect 771 -281 776 -276
rect 545 -322 550 -317
rect 701 -322 706 -317
<< pdm12contact >>
rect 76 -304 81 -299
rect 168 -304 173 -299
rect 289 -310 294 -305
rect 381 -310 386 -305
rect 577 -312 582 -307
rect 669 -312 674 -307
<< metal2 >>
rect 473 -132 490 -129
rect 473 -137 476 -132
rect 325 -168 348 -165
rect 325 -189 328 -168
rect 345 -174 348 -168
rect 765 -164 782 -161
rect 779 -169 782 -164
rect 345 -177 407 -174
rect 421 -178 483 -175
rect 236 -192 328 -189
rect 236 -214 239 -192
rect 375 -193 434 -190
rect 71 -217 239 -214
rect 71 -233 74 -217
rect 85 -226 120 -223
rect 79 -258 82 -227
rect 154 -235 158 -234
rect 154 -238 185 -235
rect 91 -244 120 -241
rect 236 -237 239 -217
rect 285 -239 288 -206
rect 375 -227 378 -193
rect 298 -232 333 -229
rect 480 -233 483 -178
rect 772 -210 834 -207
rect 762 -216 765 -210
rect 443 -237 478 -234
rect 285 -242 299 -239
rect 152 -256 177 -253
rect 304 -250 333 -247
rect 443 -243 446 -237
rect 573 -219 765 -216
rect 483 -237 528 -234
rect 374 -246 446 -243
rect 484 -248 502 -244
rect 224 -256 240 -253
rect 71 -261 82 -258
rect 71 -269 74 -261
rect 67 -272 74 -269
rect 24 -310 27 -282
rect 24 -313 44 -310
rect 63 -315 66 -273
rect 237 -269 240 -256
rect 287 -259 305 -256
rect 302 -267 305 -259
rect 302 -270 399 -267
rect 77 -287 112 -284
rect 77 -299 80 -287
rect 109 -292 112 -287
rect 137 -287 172 -284
rect 109 -295 116 -292
rect 137 -292 140 -287
rect 133 -295 140 -292
rect 169 -299 172 -287
rect 183 -315 186 -273
rect 396 -274 399 -270
rect 525 -268 528 -237
rect 573 -241 576 -219
rect 586 -234 621 -231
rect 573 -244 588 -241
rect 592 -252 621 -249
rect 658 -251 762 -248
rect 572 -262 649 -259
rect 759 -267 762 -251
rect 772 -265 775 -210
rect 821 -225 880 -222
rect 877 -259 880 -225
rect 525 -271 749 -268
rect 759 -270 772 -267
rect 205 -313 228 -310
rect 225 -339 228 -313
rect 237 -316 240 -288
rect 237 -319 257 -316
rect 276 -321 279 -279
rect 400 -278 467 -275
rect 290 -293 325 -290
rect 290 -305 293 -293
rect 322 -298 325 -293
rect 350 -293 385 -290
rect 322 -301 329 -298
rect 350 -298 353 -293
rect 346 -301 353 -298
rect 382 -305 385 -293
rect 396 -321 399 -279
rect 418 -319 441 -316
rect 438 -345 441 -319
rect 525 -318 528 -290
rect 525 -321 545 -318
rect 564 -323 567 -281
rect 746 -277 749 -271
rect 746 -280 771 -277
rect 578 -295 613 -292
rect 578 -307 581 -295
rect 610 -300 613 -295
rect 638 -295 673 -292
rect 610 -303 617 -300
rect 638 -300 641 -295
rect 634 -303 641 -300
rect 670 -307 673 -295
rect 684 -323 687 -281
rect 706 -321 729 -318
rect 726 -347 729 -321
<< m3contact >>
rect 284 -206 289 -201
rect 154 -243 159 -238
rect 434 -194 439 -189
rect 502 -249 507 -244
rect 23 -282 28 -277
rect 816 -226 821 -221
rect 236 -288 241 -283
rect 467 -279 472 -274
rect 524 -290 529 -285
<< m123contact >>
rect 122 -172 127 -167
rect 335 -178 340 -173
rect 389 -169 394 -164
rect 489 -178 494 -173
rect 433 -232 438 -227
rect 623 -180 628 -175
rect 531 -198 536 -193
rect 861 -201 866 -196
rect 122 -275 127 -270
rect 390 -261 395 -256
rect 170 -280 175 -275
rect 719 -230 724 -225
rect 843 -207 848 -202
rect 823 -264 828 -259
rect 28 -322 33 -317
rect 62 -320 67 -315
rect 182 -320 187 -315
rect 216 -322 221 -317
rect 335 -281 340 -276
rect 383 -286 388 -281
rect 241 -328 246 -323
rect 275 -326 280 -321
rect 395 -326 400 -321
rect 429 -328 434 -323
rect 623 -283 628 -278
rect 671 -288 676 -283
rect 860 -293 865 -288
rect 529 -330 534 -325
rect 563 -328 568 -323
rect 683 -328 688 -323
rect 717 -330 722 -325
<< metal3 >>
rect 380 -160 489 -157
rect 320 -164 353 -161
rect 123 -270 126 -172
rect 320 -184 323 -164
rect 350 -169 353 -164
rect 380 -169 383 -160
rect 350 -172 383 -169
rect 285 -187 323 -184
rect 285 -200 288 -187
rect 283 -201 290 -200
rect 283 -206 284 -201
rect 289 -206 290 -201
rect 283 -207 290 -206
rect 153 -238 160 -237
rect 153 -243 154 -238
rect 159 -243 160 -238
rect 153 -244 160 -243
rect 154 -260 158 -244
rect 278 -260 282 -226
rect 154 -264 282 -260
rect 22 -277 29 -276
rect 22 -282 23 -277
rect 28 -279 29 -277
rect 169 -279 170 -275
rect 28 -280 170 -279
rect 175 -280 176 -275
rect 336 -276 339 -178
rect 390 -256 393 -169
rect 486 -177 489 -160
rect 613 -170 636 -167
rect 490 -182 493 -178
rect 613 -182 616 -170
rect 633 -174 636 -170
rect 633 -177 834 -174
rect 490 -185 616 -182
rect 433 -189 440 -188
rect 433 -194 434 -189
rect 439 -190 440 -189
rect 439 -193 532 -190
rect 439 -194 440 -193
rect 433 -195 440 -194
rect 529 -196 531 -193
rect 28 -282 176 -280
rect 22 -283 29 -282
rect 235 -283 242 -282
rect 235 -288 236 -283
rect 241 -285 242 -283
rect 382 -285 383 -281
rect 241 -286 383 -285
rect 388 -286 389 -281
rect 241 -288 389 -286
rect 235 -289 242 -288
rect 434 -302 437 -232
rect 502 -243 506 -226
rect 501 -244 508 -243
rect 501 -249 502 -244
rect 507 -249 508 -244
rect 501 -250 508 -249
rect 466 -274 473 -273
rect 466 -279 467 -274
rect 472 -277 540 -274
rect 472 -279 473 -277
rect 624 -278 627 -180
rect 831 -202 834 -177
rect 831 -205 843 -202
rect 815 -221 822 -220
rect 815 -222 816 -221
rect 723 -225 816 -222
rect 724 -228 726 -225
rect 815 -226 816 -225
rect 821 -226 822 -221
rect 815 -227 822 -226
rect 813 -263 823 -260
rect 466 -280 473 -279
rect 523 -285 530 -284
rect 523 -290 524 -285
rect 529 -287 530 -285
rect 670 -287 671 -283
rect 529 -288 671 -287
rect 676 -288 677 -283
rect 813 -284 816 -263
rect 752 -287 816 -284
rect 862 -288 865 -201
rect 529 -290 677 -288
rect 523 -291 530 -290
rect 299 -305 437 -302
rect 30 -317 62 -316
rect 33 -319 62 -317
rect 187 -317 219 -316
rect 187 -319 216 -317
rect 217 -335 220 -322
rect 243 -323 275 -322
rect 246 -325 275 -323
rect 299 -335 302 -305
rect 400 -323 432 -322
rect 400 -325 429 -323
rect 531 -325 563 -324
rect 534 -327 563 -325
rect 688 -325 720 -324
rect 688 -327 717 -325
rect 217 -338 302 -335
<< m4contact >>
rect 278 -226 283 -221
rect 502 -226 507 -221
rect 540 -277 545 -272
rect 747 -288 752 -283
<< metal4 >>
rect 283 -226 502 -222
rect 545 -276 740 -273
rect 737 -285 740 -276
rect 737 -288 747 -285
<< labels >>
rlabel metal1 124 -293 124 -293 3 vdd
rlabel metal1 124 -301 124 -301 3 gnd
rlabel metal1 110 -193 110 -193 5 vdd
rlabel metal1 139 -254 139 -254 1 gnd
rlabel metal1 129 -173 129 -172 5 vdd
rlabel metal1 263 -239 269 -236 7 c1
rlabel metal1 256 -268 256 -268 1 gnd
rlabel metal1 247 -195 247 -195 5 vdd
rlabel m2contact 186 -236 190 -235 1 p0_inv
rlabel metal1 230 -232 232 -229 1 temp100
rlabel metal1 193 -173 193 -172 5 vdd
rlabel metal1 203 -254 203 -254 1 gnd
rlabel metal1 178 -210 180 -207 1 c0_inv
rlabel metal1 163 -211 165 -209 3 c0
rlabel metal1 169 -230 169 -230 1 gnd
rlabel metal1 168 -172 168 -172 5 vdd
rlabel m2contact 184 -271 185 -271 1 c0
rlabel metal2 226 -339 227 -337 1 s0
rlabel metal2 25 -312 29 -310 3 mid_s0
rlabel metal1 117 -231 128 -228 1 a0
rlabel metal1 117 -238 128 -235 1 b0
rlabel metal1 88 -237 94 -234 1 g0_inv
rlabel metal1 150 -233 155 -230 1 p0_inv
rlabel m2contact 236 -240 240 -238 1 g0_inv
rlabel metal1 337 -299 337 -299 3 vdd
rlabel metal1 337 -307 337 -307 3 gnd
rlabel metal1 323 -199 323 -199 5 vdd
rlabel metal1 352 -260 352 -260 1 gnd
rlabel metal1 342 -179 342 -178 5 vdd
rlabel metal2 238 -317 238 -317 1 mid_s1
rlabel metal2 439 -345 440 -343 8 s1
rlabel metal1 301 -243 307 -240 1 g1_inv
rlabel metal1 363 -239 368 -236 1 p1_inv
rlabel metal1 330 -237 341 -234 1 a1
rlabel metal1 330 -244 341 -241 1 b1
rlabel metal1 397 -275 399 -272 1 c1
rlabel metal1 475 -180 475 -179 5 vdd
rlabel metal1 465 -261 465 -261 1 gnd
rlabel metal1 476 -238 480 -236 7 p1_inv
rlabel metal1 477 -244 482 -242 7 p0_inv
rlabel metal1 449 -240 453 -238 3 temp101
rlabel metal1 419 -186 419 -186 5 vdd
rlabel metal1 410 -259 410 -259 1 gnd
rlabel metal1 426 -230 430 -229 1 c0
rlabel metal1 382 -229 384 -227 1 temp102
rlabel metal1 393 -157 393 -157 3 gnd
rlabel metal1 474 -167 475 -167 7 vdd
rlabel space 410 -173 413 -170 1 g0_inv
rlabel metal1 415 -131 418 -128 1 temp103
rlabel metal1 502 -132 502 -132 5 vdd
rlabel metal1 511 -205 511 -205 1 gnd
rlabel metal1 518 -176 524 -173 7 temp104
rlabel metal1 540 -132 540 -131 5 vdd
rlabel metal1 550 -213 550 -213 1 gnd
rlabel metal1 577 -191 579 -189 1 c2
rlabel m123contact 490 -176 490 -176 1 g1_inv
rlabel metal1 625 -301 625 -301 3 vdd
rlabel metal1 625 -309 625 -309 3 gnd
rlabel metal1 611 -201 611 -201 5 vdd
rlabel metal1 640 -262 640 -262 1 gnd
rlabel metal1 630 -181 630 -180 5 vdd
rlabel metal2 527 -320 528 -318 1 mid_s2
rlabel metal2 727 -347 729 -345 8 s2
rlabel metal1 618 -239 629 -236 1 a2
rlabel metal1 618 -246 629 -243 1 b2
rlabel metal1 651 -241 656 -238 1 p2_inv
rlabel metal1 760 -209 762 -207 1 g2_inv
rlabel metal1 773 -276 778 -274 1 p1_inv
rlabel metal1 837 -163 840 -160 1 temp107
rlabel metal1 775 -270 779 -268 1 p2_inv
rlabel metal1 802 -272 806 -270 1 temp105
rlabel metal1 825 -262 829 -261 1 c1
rlabel metal1 871 -261 873 -259 1 temp106
rlabel metal1 731 -208 737 -205 1 temp108
rlabel metal1 676 -223 678 -221 1 c3
rlabel metal1 705 -245 705 -245 1 gnd
rlabel metal1 715 -164 715 -163 5 vdd
rlabel metal1 744 -237 744 -237 1 gnd
rlabel metal1 753 -164 753 -164 5 vdd
rlabel metal1 780 -199 781 -199 3 vdd
rlabel metal1 862 -189 862 -189 7 gnd
rlabel metal1 845 -291 845 -291 1 gnd
rlabel metal1 836 -218 836 -218 5 vdd
rlabel metal1 790 -293 790 -293 1 gnd
rlabel metal1 780 -212 780 -211 5 vdd
rlabel m2contact 686 -279 686 -279 1 c2
rlabel m2contact 588 -244 594 -241 1 g2_inv
rlabel metal1 843 -205 846 -202 1 g1_inv
<< end >>
