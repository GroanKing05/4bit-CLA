* SPICE3 file created from bit2gen.ext - technology: scmos

.option scale=0.09u

M1000 a_223_n170# b1 vdd w_176_n176# pfet w=40 l=2
+  ad=320 pd=96 as=3180 ps=1498
M1001 p1_inv b1 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=1550 ps=880
M1002 vdd mid_s1 a_219_n261# w_235_n268# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1003 a_421_n123# temp102 vdd w_365_n109# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1004 vdd mid_s0 a_6_n255# w_22_n262# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1005 vdd g0_inv c1 w_37_n150# pfet w=20 l=2
+  ad=0 pd=0 as=260 ps=106
M1006 a_123_n204# temp100 gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1007 a_421_n151# temp102 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1008 s0 c0 mid_s0 w_61_n257# pfet w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1009 temp103 a_273_n104# vdd w_293_n89# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 g0_inv b0 vdd w_n37_n170# pfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1011 temp100 a_74_n192# vdd w_37_n150# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1012 gnd a0 a_n24_n202# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1013 gnd b0 a_n84_n281# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1014 gnd mid_s0 a_6_n255# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1015 c0 mid_s0 s0 w_61_n257# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1016 a_262_n189# c0 vdd w_250_n169# pfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1017 a_n84_n281# a0 mid_s0 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1018 temp104 temp103 vdd w_365_n109# pfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1019 temp100 a_74_n192# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1020 a_336_n171# p1_inv temp101 w_323_n177# pfet w=40 l=2
+  ad=320 pd=96 as=200 ps=90
M1021 gnd p0_inv temp101 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1022 mid_s0 a_n84_n281# a0 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1023 c1 temp100 vdd w_37_n150# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 c2 a_421_n151# vdd w_365_n109# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1025 s1 c1 a_219_n261# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1026 vdd a0 g0_inv w_n37_n170# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 gnd a1 a_189_n208# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1028 b0 a0 mid_s0 w_n95_n257# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1029 c1 a_219_n261# s1 Gnd nfet w=10 l=2
+  ad=150 pd=80 as=0 ps=0
M1030 c2 a_421_n151# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1031 a_10_n164# b0 vdd w_n37_n170# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1032 c0_inv c0 vdd w_37_n150# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1033 p0_inv b0 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1034 mid_s0 b0 a0 w_n95_n257# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1035 vdd b0 a_n84_n281# w_n55_n262# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1036 a_301_n104# g0_inv vdd w_293_n89# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1037 temp101 p1_inv gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 c0_inv c0 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1039 temp103 a_273_n104# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1040 p0_inv a0 a_10_n164# w_n37_n170# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1041 gnd a0 p0_inv Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 s1 c1 mid_s1 w_274_n263# pfet w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1043 gnd p1_inv a_273_n104# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1044 a_273_n104# p1_inv a_301_n104# w_293_n89# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1045 a_273_n104# g0_inv gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 vdd a1 g1_inv w_176_n176# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1047 a_189_n208# b1 g1_inv Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1048 c1 mid_s1 s1 w_274_n263# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 a_74_n192# c0_inv a_74_n164# w_37_n150# pfet w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1050 gnd c0_inv a_74_n192# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1051 gnd temp101 a_285_n195# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1052 temp104 g1_inv a_378_n141# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=160 ps=56
M1053 gnd mid_s1 a_219_n261# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 mid_s1 a_129_n287# a1 Gnd nfet w=10 l=2
+  ad=70 pd=34 as=50 ps=30
M1055 vdd b1 a_129_n287# w_158_n268# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1056 gnd b1 a_129_n287# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1057 a_129_n287# a1 mid_s1 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 p1_inv a1 a_223_n170# w_176_n176# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1059 gnd a1 p1_inv Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 c1 g0_inv a_123_n204# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 a_421_n151# temp104 a_421_n123# w_365_n109# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1062 gnd temp104 a_421_n151# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 a_n24_n202# b0 g0_inv Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1064 g1_inv b1 vdd w_176_n176# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 s0 c0 a_6_n255# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1066 a_74_n164# p0_inv vdd w_37_n150# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_74_n192# p0_inv gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 vdd a_262_n189# temp102 w_250_n169# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1069 a_285_n195# c0 a_262_n189# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1070 mid_s1 b1 a1 w_118_n263# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1071 a_378_n141# temp103 gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 c0 a_6_n255# s0 Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1073 vdd g1_inv temp104 w_365_n109# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 vdd temp101 a_262_n189# w_250_n169# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 b1 a1 mid_s1 w_118_n263# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1076 vdd p0_inv a_336_n171# w_323_n177# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 gnd a_262_n189# temp102 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
C0 c1 mid_s1 0.27fF
C1 c0 a_6_n255# 0.10fF
C2 g1_inv temp104 0.10fF
C3 a_273_n104# p1_inv 0.17fF
C4 gnd mid_s1 0.22fF
C5 b1 w_176_n176# 0.14fF
C6 w_118_n263# b1 0.10fF
C7 g0_inv w_n37_n170# 0.30fF
C8 g1_inv a1 0.32fF
C9 temp101 w_250_n169# 0.07fF
C10 c0 w_235_n268# 0.02fF
C11 g0_inv a_273_n104# 0.02fF
C12 vdd w_37_n150# 0.14fF
C13 b0 w_n55_n262# 0.07fF
C14 a0 w_n95_n257# 0.24fF
C15 p0_inv w_250_n169# 0.01fF
C16 temp102 a_262_n189# 0.04fF
C17 vdd g1_inv 0.04fF
C18 c0 p1_inv 0.06fF
C19 p0_inv a1 0.05fF
C20 b0 a_n24_n202# 0.01fF
C21 g0_inv c0 0.07fF
C22 b0 a0 0.71fF
C23 p0_inv a_123_n204# 0.00fF
C24 p0_inv vdd 0.09fF
C25 vdd w_293_n89# 0.09fF
C26 a_n84_n281# w_n55_n262# 0.02fF
C27 mid_s0 w_22_n262# 0.07fF
C28 b1 a_189_n208# 0.01fF
C29 temp104 w_365_n109# 0.13fF
C30 a1 mid_s1 0.40fF
C31 a0 a_n84_n281# 0.10fF
C32 c0 mid_s0 0.27fF
C33 gnd a_6_n255# 0.02fF
C34 vdd mid_s1 0.12fF
C35 a_74_n192# w_37_n150# 0.09fF
C36 p0_inv w_37_n150# 0.06fF
C37 vdd w_365_n109# 0.11fF
C38 vdd w_n55_n262# 0.11fF
C39 vdd temp103 0.84fF
C40 p0_inv g1_inv 0.06fF
C41 c0 temp102 0.00fF
C42 g1_inv w_293_n89# 0.01fF
C43 gnd p1_inv 0.20fF
C44 p0_inv a_74_n192# 0.02fF
C45 c0 b1 0.04fF
C46 g0_inv c1 0.10fF
C47 g0_inv b0 0.26fF
C48 p0_inv temp101 0.08fF
C49 c0 a_262_n189# 0.10fF
C50 g0_inv gnd 0.09fF
C51 c0 c0_inv 0.04fF
C52 a0 vdd 0.12fF
C53 mid_s0 s0 0.00fF
C54 b1 a_129_n287# 0.06fF
C55 c0 s1 0.01fF
C56 mid_s0 w_n95_n257# 0.18fF
C57 temp102 a_421_n151# 0.02fF
C58 g1_inv w_365_n109# 0.07fF
C59 b0 mid_s0 0.25fF
C60 temp103 g1_inv 0.32fF
C61 gnd mid_s0 0.22fF
C62 p1_inv a1 0.17fF
C63 vdd w_323_n177# 0.02fF
C64 vdd w_235_n268# 0.11fF
C65 temp103 w_293_n89# 0.09fF
C66 gnd temp102 0.11fF
C67 vdd p1_inv 0.56fF
C68 mid_s1 a_219_n261# 0.06fF
C69 b1 c1 0.20fF
C70 gnd b1 0.05fF
C71 a0 p0_inv 0.17fF
C72 g0_inv vdd 0.73fF
C73 gnd a_262_n189# 0.06fF
C74 c0_inv gnd 0.03fF
C75 w_274_n263# s1 0.17fF
C76 c1 s1 0.35fF
C77 c2 w_365_n109# 0.02fF
C78 c0 a_129_n287# 0.22fF
C79 temp102 a_378_n141# 0.01fF
C80 p1_inv a_285_n195# 0.01fF
C81 temp103 w_365_n109# 0.07fF
C82 temp102 w_250_n169# 0.48fF
C83 c0 s0 0.41fF
C84 vdd mid_s0 0.12fF
C85 temp102 temp104 0.24fF
C86 g1_inv p1_inv 0.05fF
C87 w_118_n263# a1 0.24fF
C88 w_158_n268# b1 0.07fF
C89 temp100 w_37_n150# 0.09fF
C90 a1 w_176_n176# 0.44fF
C91 g0_inv w_37_n150# 0.56fF
C92 b0 w_n37_n170# 0.14fF
C93 temp101 w_323_n177# 0.05fF
C94 a_262_n189# w_250_n169# 0.11fF
C95 c0 w_274_n263# 0.01fF
C96 g0_inv g1_inv 0.05fF
C97 vdd w_176_n176# 0.12fF
C98 p0_inv w_323_n177# 0.07fF
C99 p1_inv temp101 0.33fF
C100 p0_inv p1_inv 0.32fF
C101 gnd a_273_n104# 0.04fF
C102 vdd temp102 0.24fF
C103 p1_inv w_293_n89# 0.07fF
C104 b1 a1 1.02fF
C105 a_74_n192# temp100 0.04fF
C106 g0_inv a_74_n192# 0.05fF
C107 p0_inv temp100 0.00fF
C108 c0 c1 0.06fF
C109 vdd b1 0.19fF
C110 g0_inv p0_inv 0.05fF
C111 p0_inv a_336_n171# 0.01fF
C112 g0_inv w_293_n89# 0.06fF
C113 c0 gnd 0.74fF
C114 w_235_n268# a_219_n261# 0.02fF
C115 w_61_n257# mid_s0 0.10fF
C116 w_235_n268# mid_s1 0.07fF
C117 g1_inv w_176_n176# 0.04fF
C118 gnd a_421_n151# 0.04fF
C119 g1_inv temp102 0.00fF
C120 w_274_n263# c1 0.24fF
C121 g1_inv b1 0.26fF
C122 b0 w_n95_n257# 0.10fF
C123 c0 w_158_n268# 0.01fF
C124 c0 w_250_n169# 0.07fF
C125 p0_inv w_176_n176# 0.02fF
C126 vdd w_n37_n170# 0.12fF
C127 c0_inv w_37_n150# 0.12fF
C128 temp102 temp101 0.01fF
C129 p0_inv temp102 0.06fF
C130 vdd w_22_n262# 0.11fF
C131 c0_inv a_74_n192# 0.17fF
C132 c0 a1 0.01fF
C133 p0_inv b1 0.01fF
C134 g0_inv a0 0.38fF
C135 gnd c1 0.23fF
C136 p0_inv a_262_n189# 0.01fF
C137 c0 vdd 0.21fF
C138 p0_inv c0_inv 0.25fF
C139 g0_inv a_74_n164# 0.01fF
C140 b0 gnd 0.05fF
C141 w_158_n268# a_129_n287# 0.02fF
C142 a1 a_129_n287# 0.10fF
C143 temp104 a_421_n151# 0.17fF
C144 w_118_n263# mid_s1 0.18fF
C145 temp102 w_365_n109# 0.06fF
C146 b1 mid_s1 0.25fF
C147 b0 a_n84_n281# 0.06fF
C148 a0 mid_s0 0.40fF
C149 a_273_n104# g1_inv 0.07fF
C150 temp103 temp102 0.00fF
C151 p1_inv w_323_n177# 0.47fF
C152 c0 w_61_n257# 0.24fF
C153 p0_inv w_n37_n170# 0.02fF
C154 c0 w_37_n150# 0.07fF
C155 g0_inv p1_inv 0.27fF
C156 gnd w_250_n169# 0.01fF
C157 a_273_n104# w_293_n89# 0.09fF
C158 mid_s1 s1 0.00fF
C159 a1 c1 0.25fF
C160 g0_inv temp100 0.31fF
C161 p0_inv a_223_n170# 0.01fF
C162 c0 temp101 0.30fF
C163 vdd c1 0.06fF
C164 g0_inv a_10_n164# 0.01fF
C165 b0 vdd 0.19fF
C166 c0 p0_inv 0.25fF
C167 vdd gnd 1.00fF
C168 mid_s0 a_6_n255# 0.06fF
C169 w_61_n257# s0 0.17fF
C170 temp103 a_273_n104# 0.04fF
C171 p1_inv w_176_n176# 0.02fF
C172 temp102 w_323_n177# 0.01fF
C173 c0 mid_s1 0.05fF
C174 temp102 p1_inv 0.06fF
C175 c1 w_37_n150# 0.04fF
C176 a0 w_n37_n170# 0.44fF
C177 p1_inv b1 0.02fF
C178 vdd w_158_n268# 0.11fF
C179 vdd w_250_n169# 0.07fF
C180 p1_inv a_262_n189# 0.01fF
C181 temp102 a_336_n171# 0.01fF
C182 gnd g1_inv 0.06fF
C183 gnd a_74_n192# 0.04fF
C184 p0_inv c1 0.17fF
C185 vdd a1 0.12fF
C186 a_301_n104# g1_inv 0.03fF
C187 b0 p0_inv 0.02fF
C188 g0_inv c0_inv 0.12fF
C189 gnd temp101 0.02fF
C190 p0_inv gnd 0.61fF
C191 a_421_n151# c2 0.04fF
C192 c1 a_219_n261# 0.10fF
C193 a_421_n151# w_365_n109# 0.09fF
C194 gnd a_219_n261# 0.02fF
C195 w_274_n263# mid_s1 0.10fF
C196 a_6_n255# w_22_n262# 0.02fF
C197 s1 Gnd 0.43fF
C198 a_219_n261# Gnd 0.38fF
C199 a_129_n287# Gnd 0.38fF
C200 mid_s1 Gnd 1.09fF
C201 s0 Gnd 0.43fF
C202 a_6_n255# Gnd 0.38fF
C203 a_n84_n281# Gnd 0.38fF
C204 mid_s0 Gnd 1.09fF
C205 c2 Gnd 0.03fF
C206 a_421_n151# Gnd 0.18fF
C207 a_262_n189# Gnd 0.18fF
C208 temp101 Gnd 0.31fF
C209 c1 Gnd 0.07fF
C210 temp100 Gnd 0.19fF
C211 a1 Gnd 0.15fF
C212 b1 Gnd 0.07fF
C213 a_74_n192# Gnd 0.18fF
C214 gnd Gnd 3.24fF
C215 vdd Gnd 4.98fF
C216 c0_inv Gnd 0.09fF
C217 p0_inv Gnd 1.47fF
C218 c0 Gnd 0.24fF
C219 a0 Gnd 1.78fF
C220 b0 Gnd 1.19fF
C221 g0_inv Gnd 3.26fF
C222 p1_inv Gnd 2.07fF
C223 temp104 Gnd 0.28fF
C224 temp102 Gnd 0.54fF
C225 g1_inv Gnd 1.17fF
C226 a_273_n104# Gnd 0.02fF
C227 temp103 Gnd 0.49fF
C228 w_274_n263# Gnd 1.06fF
C229 w_235_n268# Gnd 0.84fF
C230 w_158_n268# Gnd 0.84fF
C231 w_118_n263# Gnd 0.42fF
C232 w_61_n257# Gnd 1.06fF
C233 w_22_n262# Gnd 0.84fF
C234 w_n55_n262# Gnd 0.84fF
C235 w_n95_n257# Gnd 1.06fF
C236 w_323_n177# Gnd 1.78fF
C237 w_250_n169# Gnd 1.43fF
C238 w_176_n176# Gnd 0.19fF
C239 w_37_n150# Gnd 1.14fF
C240 w_n37_n170# Gnd 1.09fF
C241 w_365_n109# Gnd 3.75fF
C242 w_293_n89# Gnd 2.40fF
