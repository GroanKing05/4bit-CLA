* OR Gate (inverter 2W/W)
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
* width is the universal width parameter - 10*LAMBDA
.param width = {10*LAMBDA}
.global gnd vdd

.subckt or in_1 in_2 out width
    * NOR gate
    MP1 temp1 in_1 vdd vdd CMOSP W={(2*width)} L={2*LAMBDA}
    + AS={5*(2*width)*LAMBDA} PS={10*LAMBDA+2*(2*width)} AD={5*(2*width)*LAMBDA} PD={10*LAMBDA+2*(2*width)}
    MP2 out1 in_2 temp1 vdd CMOSP W={(2*width)} L={2*LAMBDA}
    + AS={5*(2*width)*LAMBDA} PS={10*LAMBDA+2*(2*width)} AD={5*(2*width)*LAMBDA} PD={10*LAMBDA+2*(2*width)}
    MN1 out1 in_1 gnd gnd CMOSN W={(2*width)} L={2*LAMBDA}
    + AS={5*(2*width)*LAMBDA} PS={10*LAMBDA+2*(2*width)} AD={5*(2*width)*LAMBDA} PD={10*LAMBDA+2*(2*width)}
    MN2 out1 in_2 gnd gnd CMOSN W={(2*width)} L={2*LAMBDA}
    + AS={5*(2*width)*LAMBDA} PS={10*LAMBDA+2*(2*width)} AD={5*(2*width)*LAMBDA} PD={10*LAMBDA+2*(2*width)}

    * Inverter
    MP3 out out1 vdd vdd CMOSP W={(2*width)} L={2*LAMBDA}
    + AS={5*(2*width)*LAMBDA} PS={10*LAMBDA+2*(2*width)} AD={5*(2*width)*LAMBDA} PD={10*LAMBDA+2*(2*width)}
    MN3 out out1 gnd gnd CMOSN W={(width)} L={2*LAMBDA}
    + AS={5*(width)*LAMBDA} PS={10*LAMBDA+2*(width)} AD={5*(width)*LAMBDA} PD={10*LAMBDA+2*(width)}
.ends or

Vdd vdd gnd 'SUPPLY'
Va a gnd pulse 0 1.8 0 0.01ns 0.01ns 10ns 20ns
Vb b gnd pulse 0 1.8 0 0.01ns 0.01ns 20ns 40ns

X1 a b z width or

.tran 100p 50n

.control
set hcopypscolor = 1
set color0=white
set color1=black

run

set curplottitle="2023112005_OR"
plot v(a)+2, v(b)+4, v(z)
.endc