magic
tech scmos
timestamp 1731406662
<< nwell >>
rect -94 -167 -61 -135
rect -54 -156 -22 -130
rect 23 -156 55 -130
rect 62 -167 95 -135
<< ntransistor >>
rect -83 -128 -81 -118
rect -74 -128 -72 -118
rect 73 -128 75 -118
rect 82 -128 84 -118
rect -16 -144 -6 -142
rect 7 -144 17 -142
<< ptransistor >>
rect -83 -161 -81 -141
rect -74 -161 -72 -141
rect -48 -144 -28 -142
rect 29 -144 49 -142
rect 73 -161 75 -141
rect 82 -161 84 -141
<< ndiffusion >>
rect -88 -124 -83 -118
rect -84 -128 -83 -124
rect -81 -124 -74 -118
rect -81 -128 -79 -124
rect -75 -128 -74 -124
rect -72 -122 -71 -118
rect -72 -128 -67 -122
rect 72 -122 73 -118
rect 68 -128 73 -122
rect 75 -124 82 -118
rect 75 -128 76 -124
rect 80 -128 82 -124
rect 84 -124 89 -118
rect 84 -128 85 -124
rect -12 -141 -6 -137
rect -16 -142 -6 -141
rect 7 -141 13 -137
rect 7 -142 17 -141
rect -16 -145 -6 -144
rect -16 -149 -10 -145
rect 7 -145 17 -144
rect 11 -149 17 -145
<< pdiffusion >>
rect -48 -141 -32 -137
rect -84 -145 -83 -141
rect -88 -161 -83 -145
rect -81 -143 -74 -141
rect -81 -147 -79 -143
rect -75 -147 -74 -143
rect -81 -161 -74 -147
rect -72 -157 -67 -141
rect -48 -142 -28 -141
rect 33 -141 49 -137
rect 29 -142 49 -141
rect -48 -145 -28 -144
rect -43 -150 -28 -145
rect 29 -145 49 -144
rect 29 -150 44 -145
rect -72 -161 -71 -157
rect 68 -157 73 -141
rect 72 -161 73 -157
rect 75 -143 82 -141
rect 75 -147 76 -143
rect 80 -147 82 -143
rect 75 -161 82 -147
rect 84 -145 85 -141
rect 84 -161 89 -145
<< ndcontact >>
rect -88 -128 -84 -124
rect -79 -128 -75 -124
rect -71 -122 -67 -118
rect 68 -122 72 -118
rect 76 -128 80 -124
rect 85 -128 89 -124
rect -16 -141 -12 -137
rect 13 -141 17 -137
rect -10 -149 -6 -145
rect 7 -149 11 -145
<< pdcontact >>
rect -32 -141 -28 -137
rect -88 -145 -84 -141
rect -79 -147 -75 -143
rect 29 -141 33 -137
rect -71 -161 -67 -157
rect 68 -161 72 -157
rect 76 -147 80 -143
rect 85 -145 89 -141
<< polysilicon >>
rect -83 -112 -81 -111
rect 82 -112 84 -111
rect -83 -116 -82 -112
rect -83 -118 -81 -116
rect -74 -118 -72 -115
rect 73 -118 75 -115
rect 83 -116 84 -112
rect 82 -118 84 -116
rect -83 -132 -81 -128
rect -83 -141 -81 -135
rect -74 -141 -72 -128
rect 73 -141 75 -128
rect 82 -132 84 -128
rect 82 -141 84 -135
rect -52 -144 -48 -142
rect -28 -144 -16 -142
rect -6 -144 -2 -142
rect 3 -144 7 -142
rect 17 -144 29 -142
rect 49 -144 53 -142
rect -83 -173 -81 -161
rect -74 -164 -72 -161
rect 73 -164 75 -161
rect 82 -173 84 -161
<< polycontact >>
rect -82 -116 -78 -112
rect 79 -116 83 -112
rect -72 -134 -68 -130
rect 69 -134 73 -130
rect -21 -148 -17 -144
rect 18 -148 22 -144
rect -81 -172 -77 -168
rect 78 -172 82 -168
<< metal1 >>
rect -78 -115 -61 -112
rect -64 -118 -61 -115
rect -67 -120 -61 -118
rect 62 -115 79 -112
rect 62 -118 65 -115
rect 62 -120 68 -118
rect -67 -121 -48 -120
rect -64 -123 -48 -121
rect -87 -131 -84 -128
rect -91 -132 -84 -131
rect -96 -134 -84 -132
rect -87 -141 -84 -134
rect -51 -126 -48 -123
rect 49 -121 68 -120
rect 49 -123 65 -121
rect 49 -126 52 -123
rect -79 -135 -76 -128
rect -51 -129 -18 -126
rect -68 -133 -62 -130
rect -21 -137 -18 -129
rect 19 -129 52 -126
rect 19 -137 22 -129
rect 63 -133 69 -130
rect 77 -135 80 -128
rect 85 -131 88 -128
rect 85 -132 92 -131
rect 85 -134 97 -132
rect -79 -143 -76 -140
rect -28 -140 -16 -137
rect 17 -140 29 -137
rect 77 -143 80 -140
rect -21 -158 -18 -148
rect -6 -149 7 -146
rect -3 -157 4 -154
rect 19 -158 22 -148
rect 85 -141 88 -134
rect -67 -161 -18 -158
rect 19 -161 68 -158
rect -58 -168 -55 -161
rect -51 -168 -44 -167
rect 56 -168 59 -161
rect -77 -169 -44 -168
rect -77 -171 -50 -169
rect -51 -174 -50 -171
rect -45 -174 -44 -169
rect 47 -171 78 -168
rect -61 -183 -58 -181
rect 47 -183 50 -171
rect 59 -183 62 -181
<< m2contact >>
rect -80 -140 -75 -135
rect 76 -140 81 -135
rect -8 -158 -3 -153
rect 4 -158 9 -153
rect -62 -181 -57 -176
rect 58 -181 63 -176
<< pdm12contact >>
rect -48 -150 -43 -145
rect 44 -150 49 -145
<< metal2 >>
rect -103 -136 -100 -110
rect -103 -139 -80 -136
rect -61 -176 -58 -134
rect -47 -162 -44 -150
rect -15 -157 -8 -154
rect -15 -162 -12 -157
rect 9 -157 16 -154
rect -47 -165 -12 -162
rect 13 -162 16 -157
rect 45 -162 48 -150
rect 13 -165 48 -162
rect 59 -176 62 -134
rect 81 -139 101 -136
rect 98 -167 101 -139
<< m3contact >>
rect 97 -172 102 -167
<< m123contact >>
rect -96 -132 -91 -127
rect -62 -134 -57 -129
rect 58 -134 63 -129
rect 92 -132 97 -127
rect -50 -174 -45 -169
<< metal3 >>
rect -91 -132 -62 -130
rect -94 -133 -62 -132
rect 63 -132 92 -130
rect 63 -133 95 -132
rect 96 -167 103 -166
rect -51 -169 97 -167
rect -51 -174 -50 -169
rect -45 -170 97 -169
rect -45 -174 -44 -170
rect 96 -172 97 -170
rect 102 -172 103 -167
rect 96 -173 103 -172
<< labels >>
rlabel metal1 48 -182 48 -182 1 in1
rlabel metal1 60 -182 60 -182 1 in2
rlabel metal1 1 -156 1 -156 7 vdd
rlabel metal1 1 -148 1 -148 7 gnd
rlabel metal2 98 -138 99 -138 7 mid_sumbit
rlabel metal1 -61 -183 -59 -180 1 carry_in
rlabel metal2 -102 -111 -102 -111 3 sum_bit
<< end >>
