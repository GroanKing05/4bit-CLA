magic
tech scmos
timestamp 1731350567
<< nwell >>
rect -1 62 33 68
rect -1 36 55 62
rect 30 30 55 36
<< ntransistor >>
rect 10 4 12 24
rect 20 4 22 24
rect 41 14 43 24
<< ptransistor >>
rect 10 42 12 62
rect 20 42 22 62
rect 41 36 43 56
<< ndiffusion >>
rect 5 8 10 24
rect 9 4 10 8
rect 12 4 20 24
rect 22 20 23 24
rect 22 4 27 20
rect 36 18 41 24
rect 40 14 41 18
rect 43 20 44 24
rect 43 14 48 20
<< pdiffusion >>
rect 9 58 10 62
rect 5 42 10 58
rect 12 46 20 62
rect 12 42 14 46
rect 18 42 20 46
rect 22 58 23 62
rect 22 42 27 58
rect 40 52 41 56
rect 36 36 41 52
rect 43 40 48 56
rect 43 36 44 40
<< ndcontact >>
rect 5 4 9 8
rect 23 20 27 24
rect 36 14 40 18
rect 44 20 48 24
<< pdcontact >>
rect 5 58 9 62
rect 14 42 18 46
rect 23 58 27 62
rect 36 52 40 56
rect 44 36 48 40
<< polysilicon >>
rect 10 62 12 66
rect 20 62 22 66
rect 41 56 43 60
rect 10 24 12 42
rect 20 24 22 42
rect 41 24 43 36
rect 41 10 43 14
rect 10 0 12 4
rect 20 0 22 4
<< polycontact >>
rect 6 31 10 35
rect 16 25 20 29
rect 37 25 41 29
<< metal1 >>
rect -1 69 39 72
rect 5 62 8 69
rect 23 62 27 69
rect 36 56 39 69
rect 15 41 18 42
rect 15 38 27 41
rect -1 32 6 35
rect 24 29 27 38
rect 45 29 48 36
rect -1 25 16 28
rect 24 26 37 29
rect 24 24 27 26
rect 45 26 52 29
rect 45 24 48 26
rect 5 -1 8 4
rect 36 -1 39 14
rect -1 -4 39 -1
<< labels >>
rlabel metal1 11 70 11 70 5 vdd
rlabel metal1 2 33 3 34 1 in1
rlabel metal1 2 26 2 27 1 in2
rlabel metal1 20 -3 20 -3 1 gnd
rlabel metal1 47 28 47 28 1 out
<< end >>
