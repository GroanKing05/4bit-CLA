magic
tech scmos
timestamp 1731468930
<< nwell >>
rect -885 -526 -743 -494
rect -290 -551 -258 -532
rect -290 -557 -236 -551
rect -887 -613 -745 -581
rect -288 -585 -236 -557
rect -218 -567 -141 -545
rect 803 -547 945 -515
rect 954 -548 979 -516
rect -218 -577 -123 -567
rect -586 -606 -552 -586
rect -620 -638 -552 -606
rect -546 -608 -488 -586
rect -546 -618 -439 -608
rect -373 -612 -339 -592
rect -311 -605 -277 -599
rect -522 -638 -439 -618
rect -494 -640 -439 -638
rect -407 -644 -339 -612
rect -333 -631 -277 -605
rect -333 -637 -308 -631
rect -260 -645 -226 -593
rect -175 -597 -123 -577
rect -147 -599 -123 -597
rect -85 -614 -51 -594
rect -20 -599 57 -577
rect 97 -583 129 -564
rect -119 -646 -51 -614
rect -38 -609 57 -599
rect 75 -589 129 -583
rect -38 -629 14 -609
rect 75 -617 127 -589
rect 276 -618 310 -598
rect -38 -631 -14 -629
rect -891 -704 -749 -672
rect 65 -677 99 -625
rect 116 -637 150 -631
rect 116 -663 172 -637
rect 242 -650 310 -618
rect 326 -601 360 -596
rect 326 -607 397 -601
rect 326 -633 419 -607
rect 453 -621 487 -601
rect 453 -623 521 -621
rect 326 -648 360 -633
rect 394 -639 419 -633
rect 434 -627 521 -623
rect 434 -653 542 -627
rect 434 -655 459 -653
rect 518 -659 542 -653
rect 553 -633 587 -611
rect 553 -663 606 -633
rect 147 -669 172 -663
rect 581 -665 606 -663
rect 612 -665 646 -633
rect 801 -634 943 -602
rect 951 -635 976 -603
rect -678 -725 -645 -693
rect -638 -730 -606 -704
rect -561 -730 -529 -704
rect -522 -725 -489 -693
rect -465 -731 -432 -699
rect -425 -736 -393 -710
rect -348 -736 -316 -710
rect -309 -731 -276 -699
rect -177 -733 -144 -701
rect -137 -738 -105 -712
rect -60 -738 -28 -712
rect -21 -733 12 -701
rect 184 -737 217 -705
rect 224 -742 256 -716
rect 301 -742 333 -716
rect 340 -737 373 -705
rect -894 -791 -752 -759
rect 425 -776 457 -708
rect 534 -737 586 -703
rect 797 -726 939 -694
rect 950 -727 975 -695
rect 794 -812 936 -780
rect 951 -813 976 -781
rect -893 -888 -751 -856
rect 795 -909 937 -877
rect 949 -910 974 -878
rect -895 -978 -753 -946
rect -896 -1068 -754 -1036
rect -897 -1160 -755 -1128
rect -895 -1256 -753 -1224
<< ntransistor >>
rect -874 -552 -872 -532
rect -850 -552 -848 -532
rect -824 -546 -822 -536
rect -806 -552 -804 -532
rect -797 -552 -795 -532
rect -781 -552 -779 -532
rect -772 -552 -770 -532
rect -756 -546 -754 -536
rect -306 -546 -296 -544
rect -310 -564 -300 -562
rect -310 -574 -300 -572
rect -876 -639 -874 -619
rect -852 -639 -850 -619
rect -826 -633 -824 -623
rect -808 -639 -806 -619
rect -799 -639 -797 -619
rect -783 -639 -781 -619
rect -774 -639 -772 -619
rect -758 -633 -756 -623
rect -535 -634 -533 -624
rect -609 -670 -607 -650
rect -599 -670 -597 -650
rect -575 -660 -573 -650
rect -565 -660 -563 -650
rect -511 -660 -509 -650
rect -501 -660 -499 -650
rect -483 -656 -481 -646
rect -462 -672 -460 -652
rect -452 -672 -450 -652
rect -207 -609 -205 -589
rect -197 -609 -195 -589
rect 814 -573 816 -553
rect 135 -578 145 -576
rect 838 -573 840 -553
rect -164 -619 -162 -609
rect -154 -619 -152 -609
rect -136 -615 -134 -605
rect -321 -653 -319 -643
rect -396 -676 -394 -656
rect -386 -676 -384 -656
rect -362 -666 -360 -656
rect -352 -666 -350 -656
rect -300 -663 -298 -643
rect -290 -663 -288 -643
rect 864 -567 866 -557
rect 882 -573 884 -553
rect 891 -573 893 -553
rect 907 -573 909 -553
rect 916 -573 918 -553
rect 932 -567 934 -557
rect 965 -564 967 -554
rect 139 -596 149 -594
rect 139 -606 149 -604
rect -249 -667 -247 -657
rect -239 -667 -237 -657
rect -27 -647 -25 -637
rect 34 -641 36 -621
rect 44 -641 46 -621
rect -9 -651 -7 -641
rect 1 -651 3 -641
rect -108 -678 -106 -658
rect -98 -678 -96 -658
rect -74 -668 -72 -658
rect -64 -668 -62 -658
rect -880 -730 -878 -710
rect -856 -730 -854 -710
rect -830 -724 -828 -714
rect -812 -730 -810 -710
rect -803 -730 -801 -710
rect -787 -730 -785 -710
rect -778 -730 -776 -710
rect -762 -724 -760 -714
rect -600 -718 -590 -716
rect -577 -718 -567 -716
rect -387 -724 -377 -722
rect -364 -724 -354 -722
rect -667 -742 -665 -732
rect -658 -742 -656 -732
rect -511 -742 -509 -732
rect -502 -742 -500 -732
rect 76 -699 78 -689
rect 86 -699 88 -689
rect 127 -695 129 -675
rect 137 -695 139 -675
rect 158 -685 160 -675
rect 253 -682 255 -662
rect 263 -682 265 -662
rect 287 -672 289 -662
rect 297 -672 299 -662
rect 337 -670 339 -660
rect 347 -670 349 -660
rect 374 -665 376 -645
rect 384 -665 386 -645
rect 405 -655 407 -645
rect 446 -671 448 -661
rect 464 -675 466 -665
rect 474 -675 476 -665
rect 498 -685 500 -665
rect 508 -685 510 -665
rect 529 -675 531 -665
rect 564 -685 566 -675
rect 574 -685 576 -675
rect 592 -681 594 -671
rect 812 -660 814 -640
rect 836 -660 838 -640
rect 862 -654 864 -644
rect 880 -660 882 -640
rect 889 -660 891 -640
rect 905 -660 907 -640
rect 914 -660 916 -640
rect 930 -654 932 -644
rect 962 -651 964 -641
rect 623 -697 625 -677
rect 633 -697 635 -677
rect -99 -726 -89 -724
rect -76 -726 -66 -724
rect -454 -748 -452 -738
rect -445 -748 -443 -738
rect -298 -748 -296 -738
rect -289 -748 -287 -738
rect 262 -730 272 -728
rect 285 -730 295 -728
rect -166 -750 -164 -740
rect -157 -750 -155 -740
rect -10 -750 -8 -740
rect -1 -750 1 -740
rect 598 -716 608 -714
rect 469 -721 489 -719
rect 598 -726 608 -724
rect 469 -731 489 -729
rect 195 -754 197 -744
rect 204 -754 206 -744
rect 351 -754 353 -744
rect 360 -754 362 -744
rect 808 -752 810 -732
rect 469 -755 489 -753
rect 832 -752 834 -732
rect 469 -765 489 -763
rect 858 -746 860 -736
rect 876 -752 878 -732
rect 885 -752 887 -732
rect 901 -752 903 -732
rect 910 -752 912 -732
rect 926 -746 928 -736
rect 961 -743 963 -733
rect -883 -817 -881 -797
rect -859 -817 -857 -797
rect -833 -811 -831 -801
rect -815 -817 -813 -797
rect -806 -817 -804 -797
rect -790 -817 -788 -797
rect -781 -817 -779 -797
rect -765 -811 -763 -801
rect 805 -838 807 -818
rect 829 -838 831 -818
rect 855 -832 857 -822
rect 873 -838 875 -818
rect 882 -838 884 -818
rect 898 -838 900 -818
rect 907 -838 909 -818
rect 923 -832 925 -822
rect 962 -829 964 -819
rect -882 -914 -880 -894
rect -858 -914 -856 -894
rect -832 -908 -830 -898
rect -814 -914 -812 -894
rect -805 -914 -803 -894
rect -789 -914 -787 -894
rect -780 -914 -778 -894
rect -764 -908 -762 -898
rect 806 -935 808 -915
rect 830 -935 832 -915
rect 856 -929 858 -919
rect 874 -935 876 -915
rect 883 -935 885 -915
rect 899 -935 901 -915
rect 908 -935 910 -915
rect 924 -929 926 -919
rect 960 -926 962 -916
rect -884 -1004 -882 -984
rect -860 -1004 -858 -984
rect -834 -998 -832 -988
rect -816 -1004 -814 -984
rect -807 -1004 -805 -984
rect -791 -1004 -789 -984
rect -782 -1004 -780 -984
rect -766 -998 -764 -988
rect -885 -1094 -883 -1074
rect -861 -1094 -859 -1074
rect -835 -1088 -833 -1078
rect -817 -1094 -815 -1074
rect -808 -1094 -806 -1074
rect -792 -1094 -790 -1074
rect -783 -1094 -781 -1074
rect -767 -1088 -765 -1078
rect -886 -1186 -884 -1166
rect -862 -1186 -860 -1166
rect -836 -1180 -834 -1170
rect -818 -1186 -816 -1166
rect -809 -1186 -807 -1166
rect -793 -1186 -791 -1166
rect -784 -1186 -782 -1166
rect -768 -1180 -766 -1170
rect -884 -1282 -882 -1262
rect -860 -1282 -858 -1262
rect -834 -1276 -832 -1266
rect -816 -1282 -814 -1262
rect -807 -1282 -805 -1262
rect -791 -1282 -789 -1262
rect -782 -1282 -780 -1262
rect -766 -1276 -764 -1266
<< ptransistor >>
rect -874 -520 -872 -500
rect -866 -520 -864 -500
rect -850 -520 -848 -500
rect -842 -520 -840 -500
rect -824 -520 -822 -500
rect -806 -520 -804 -500
rect -781 -520 -779 -500
rect -756 -520 -754 -500
rect 814 -541 816 -521
rect 822 -541 824 -521
rect 838 -541 840 -521
rect 846 -541 848 -521
rect 864 -541 866 -521
rect 882 -541 884 -521
rect 907 -541 909 -521
rect 932 -541 934 -521
rect -284 -546 -264 -544
rect -282 -564 -242 -562
rect -207 -571 -205 -551
rect -197 -571 -195 -551
rect -282 -574 -242 -572
rect -876 -607 -874 -587
rect -868 -607 -866 -587
rect -852 -607 -850 -587
rect -844 -607 -842 -587
rect -826 -607 -824 -587
rect -808 -607 -806 -587
rect -783 -607 -781 -587
rect -758 -607 -756 -587
rect -609 -632 -607 -612
rect -599 -632 -597 -612
rect -575 -632 -573 -592
rect -565 -632 -563 -592
rect -535 -612 -533 -592
rect -511 -632 -509 -592
rect -501 -632 -499 -592
rect -483 -634 -481 -614
rect -462 -634 -460 -614
rect -452 -634 -450 -614
rect -396 -638 -394 -618
rect -386 -638 -384 -618
rect -362 -638 -360 -598
rect -352 -638 -350 -598
rect -321 -631 -319 -611
rect -300 -625 -298 -605
rect -290 -625 -288 -605
rect -249 -639 -247 -599
rect -239 -639 -237 -599
rect -164 -591 -162 -551
rect -154 -591 -152 -551
rect -136 -593 -134 -573
rect 103 -578 123 -576
rect -108 -640 -106 -620
rect -98 -640 -96 -620
rect -74 -640 -72 -600
rect -64 -640 -62 -600
rect -27 -625 -25 -605
rect -9 -623 -7 -583
rect 1 -623 3 -583
rect 34 -603 36 -583
rect 44 -603 46 -583
rect 965 -542 967 -522
rect 81 -596 121 -594
rect 81 -606 121 -604
rect -880 -698 -878 -678
rect -872 -698 -870 -678
rect -856 -698 -854 -678
rect -848 -698 -846 -678
rect -830 -698 -828 -678
rect -812 -698 -810 -678
rect -787 -698 -785 -678
rect -762 -698 -760 -678
rect 76 -671 78 -631
rect 86 -671 88 -631
rect 127 -657 129 -637
rect 137 -657 139 -637
rect 158 -663 160 -643
rect 253 -644 255 -624
rect 263 -644 265 -624
rect 287 -644 289 -604
rect 297 -644 299 -604
rect 337 -642 339 -602
rect 347 -642 349 -602
rect 374 -627 376 -607
rect 384 -627 386 -607
rect 405 -633 407 -613
rect -667 -719 -665 -699
rect -658 -719 -656 -699
rect -632 -718 -612 -716
rect -555 -718 -535 -716
rect -511 -719 -509 -699
rect -502 -719 -500 -699
rect -454 -725 -452 -705
rect -445 -725 -443 -705
rect -419 -724 -399 -722
rect -342 -724 -322 -722
rect -298 -725 -296 -705
rect -289 -725 -287 -705
rect 446 -649 448 -629
rect 464 -647 466 -607
rect 474 -647 476 -607
rect 498 -647 500 -627
rect 508 -647 510 -627
rect 529 -653 531 -633
rect 564 -657 566 -617
rect 574 -657 576 -617
rect 812 -628 814 -608
rect 820 -628 822 -608
rect 836 -628 838 -608
rect 844 -628 846 -608
rect 862 -628 864 -608
rect 880 -628 882 -608
rect 905 -628 907 -608
rect 930 -628 932 -608
rect 592 -659 594 -639
rect 623 -659 625 -639
rect 633 -659 635 -639
rect 962 -629 964 -609
rect -166 -727 -164 -707
rect -157 -727 -155 -707
rect -131 -726 -111 -724
rect -54 -726 -34 -724
rect -10 -727 -8 -707
rect -1 -727 1 -707
rect 195 -731 197 -711
rect 204 -731 206 -711
rect 230 -730 250 -728
rect 307 -730 327 -728
rect 351 -731 353 -711
rect 360 -731 362 -711
rect 540 -716 580 -714
rect 431 -721 451 -719
rect 808 -720 810 -700
rect 816 -720 818 -700
rect 832 -720 834 -700
rect 840 -720 842 -700
rect 858 -720 860 -700
rect 876 -720 878 -700
rect 901 -720 903 -700
rect 926 -720 928 -700
rect 540 -726 580 -724
rect 431 -731 451 -729
rect 431 -755 451 -753
rect 431 -765 451 -763
rect 961 -721 963 -701
rect -883 -785 -881 -765
rect -875 -785 -873 -765
rect -859 -785 -857 -765
rect -851 -785 -849 -765
rect -833 -785 -831 -765
rect -815 -785 -813 -765
rect -790 -785 -788 -765
rect -765 -785 -763 -765
rect 805 -806 807 -786
rect 813 -806 815 -786
rect 829 -806 831 -786
rect 837 -806 839 -786
rect 855 -806 857 -786
rect 873 -806 875 -786
rect 898 -806 900 -786
rect 923 -806 925 -786
rect 962 -807 964 -787
rect -882 -882 -880 -862
rect -874 -882 -872 -862
rect -858 -882 -856 -862
rect -850 -882 -848 -862
rect -832 -882 -830 -862
rect -814 -882 -812 -862
rect -789 -882 -787 -862
rect -764 -882 -762 -862
rect 806 -903 808 -883
rect 814 -903 816 -883
rect 830 -903 832 -883
rect 838 -903 840 -883
rect 856 -903 858 -883
rect 874 -903 876 -883
rect 899 -903 901 -883
rect 924 -903 926 -883
rect 960 -904 962 -884
rect -884 -972 -882 -952
rect -876 -972 -874 -952
rect -860 -972 -858 -952
rect -852 -972 -850 -952
rect -834 -972 -832 -952
rect -816 -972 -814 -952
rect -791 -972 -789 -952
rect -766 -972 -764 -952
rect -885 -1062 -883 -1042
rect -877 -1062 -875 -1042
rect -861 -1062 -859 -1042
rect -853 -1062 -851 -1042
rect -835 -1062 -833 -1042
rect -817 -1062 -815 -1042
rect -792 -1062 -790 -1042
rect -767 -1062 -765 -1042
rect -886 -1154 -884 -1134
rect -878 -1154 -876 -1134
rect -862 -1154 -860 -1134
rect -854 -1154 -852 -1134
rect -836 -1154 -834 -1134
rect -818 -1154 -816 -1134
rect -793 -1154 -791 -1134
rect -768 -1154 -766 -1134
rect -884 -1250 -882 -1230
rect -876 -1250 -874 -1230
rect -860 -1250 -858 -1230
rect -852 -1250 -850 -1230
rect -834 -1250 -832 -1230
rect -816 -1250 -814 -1230
rect -791 -1250 -789 -1230
rect -766 -1250 -764 -1230
<< ndiffusion >>
rect -879 -548 -874 -532
rect -875 -552 -874 -548
rect -872 -536 -871 -532
rect -872 -552 -867 -536
rect -855 -548 -850 -532
rect -851 -552 -850 -548
rect -848 -536 -847 -532
rect -848 -552 -843 -536
rect -829 -542 -824 -536
rect -825 -546 -824 -542
rect -822 -540 -821 -536
rect -822 -546 -817 -540
rect -811 -548 -806 -532
rect -807 -552 -806 -548
rect -804 -552 -797 -532
rect -795 -536 -794 -532
rect -795 -552 -790 -536
rect -786 -548 -781 -532
rect -782 -552 -781 -548
rect -779 -552 -772 -532
rect -770 -536 -769 -532
rect -770 -552 -765 -536
rect -761 -542 -756 -536
rect -757 -546 -756 -542
rect -754 -540 -753 -536
rect -754 -546 -749 -540
rect -306 -543 -300 -539
rect -306 -544 -296 -543
rect -306 -547 -296 -546
rect -302 -551 -296 -547
rect -306 -561 -300 -557
rect -310 -562 -300 -561
rect -310 -566 -300 -564
rect -310 -570 -304 -566
rect -310 -572 -300 -570
rect -310 -575 -300 -574
rect -306 -579 -300 -575
rect -881 -635 -876 -619
rect -877 -639 -876 -635
rect -874 -623 -873 -619
rect -874 -639 -869 -623
rect -857 -635 -852 -619
rect -853 -639 -852 -635
rect -850 -623 -849 -619
rect -850 -639 -845 -623
rect -831 -629 -826 -623
rect -827 -633 -826 -629
rect -824 -627 -823 -623
rect -824 -633 -819 -627
rect -813 -635 -808 -619
rect -809 -639 -808 -635
rect -806 -639 -799 -619
rect -797 -623 -796 -619
rect -797 -639 -792 -623
rect -788 -635 -783 -619
rect -784 -639 -783 -635
rect -781 -639 -774 -619
rect -772 -623 -771 -619
rect -772 -639 -767 -623
rect -763 -629 -758 -623
rect -759 -633 -758 -629
rect -756 -627 -755 -623
rect -756 -633 -751 -627
rect -540 -630 -535 -624
rect -536 -634 -535 -630
rect -533 -628 -532 -624
rect -533 -634 -528 -628
rect -610 -654 -609 -650
rect -614 -670 -609 -654
rect -607 -670 -599 -650
rect -597 -666 -592 -650
rect -580 -656 -575 -650
rect -576 -660 -575 -656
rect -573 -654 -571 -650
rect -567 -654 -565 -650
rect -573 -660 -565 -654
rect -563 -656 -558 -650
rect -563 -660 -562 -656
rect -516 -656 -511 -650
rect -512 -660 -511 -656
rect -509 -654 -507 -650
rect -503 -654 -501 -650
rect -509 -660 -501 -654
rect -499 -656 -494 -650
rect -488 -652 -483 -646
rect -484 -656 -483 -652
rect -481 -650 -480 -646
rect -481 -656 -476 -650
rect -499 -660 -498 -656
rect -597 -670 -596 -666
rect -467 -668 -462 -652
rect -463 -672 -462 -668
rect -460 -672 -452 -652
rect -450 -656 -449 -652
rect -212 -605 -207 -589
rect -208 -609 -207 -605
rect -205 -609 -197 -589
rect -195 -593 -194 -589
rect 809 -569 814 -553
rect -195 -609 -190 -593
rect 139 -575 145 -571
rect 813 -573 814 -569
rect 816 -557 817 -553
rect 816 -573 821 -557
rect 135 -576 145 -575
rect 135 -579 145 -578
rect 135 -583 141 -579
rect 833 -569 838 -553
rect 837 -573 838 -569
rect 840 -557 841 -553
rect 840 -573 845 -557
rect -169 -615 -164 -609
rect -165 -619 -164 -615
rect -162 -613 -160 -609
rect -156 -613 -154 -609
rect -162 -619 -154 -613
rect -152 -615 -147 -609
rect -141 -611 -136 -605
rect -137 -615 -136 -611
rect -134 -609 -133 -605
rect -134 -615 -129 -609
rect -152 -619 -151 -615
rect -322 -647 -321 -643
rect -326 -653 -321 -647
rect -319 -649 -314 -643
rect -319 -653 -318 -649
rect -301 -647 -300 -643
rect -450 -672 -445 -656
rect -397 -660 -396 -656
rect -401 -676 -396 -660
rect -394 -676 -386 -656
rect -384 -672 -379 -656
rect -367 -662 -362 -656
rect -363 -666 -362 -662
rect -360 -660 -358 -656
rect -354 -660 -352 -656
rect -360 -666 -352 -660
rect -350 -662 -345 -656
rect -350 -666 -349 -662
rect -305 -663 -300 -647
rect -298 -663 -290 -643
rect -288 -659 -283 -643
rect 859 -563 864 -557
rect 863 -567 864 -563
rect 866 -561 867 -557
rect 866 -567 871 -561
rect 877 -569 882 -553
rect 881 -573 882 -569
rect 884 -573 891 -553
rect 893 -557 894 -553
rect 893 -573 898 -557
rect 902 -569 907 -553
rect 906 -573 907 -569
rect 909 -573 916 -553
rect 918 -557 919 -553
rect 918 -573 923 -557
rect 927 -563 932 -557
rect 931 -567 932 -563
rect 934 -561 935 -557
rect 934 -567 939 -561
rect 960 -560 965 -554
rect 964 -564 965 -560
rect 967 -558 968 -554
rect 967 -564 972 -558
rect 139 -593 145 -589
rect 139 -594 149 -593
rect 139 -598 149 -596
rect 143 -602 149 -598
rect 139 -604 149 -602
rect 139 -607 149 -606
rect 139 -611 145 -607
rect -288 -663 -287 -659
rect -254 -663 -249 -657
rect -250 -667 -249 -663
rect -247 -661 -245 -657
rect -241 -661 -239 -657
rect -247 -667 -239 -661
rect -237 -663 -232 -657
rect -28 -641 -27 -637
rect -32 -647 -27 -641
rect -25 -643 -20 -637
rect 33 -625 34 -621
rect 29 -641 34 -625
rect 36 -641 44 -621
rect 46 -637 51 -621
rect 46 -641 47 -637
rect -25 -647 -24 -643
rect -14 -647 -9 -641
rect -10 -651 -9 -647
rect -7 -645 -5 -641
rect -1 -645 1 -641
rect -7 -651 1 -645
rect 3 -647 8 -641
rect 3 -651 4 -647
rect -237 -667 -236 -663
rect -109 -662 -108 -658
rect -384 -676 -383 -672
rect -113 -678 -108 -662
rect -106 -678 -98 -658
rect -96 -674 -91 -658
rect -79 -664 -74 -658
rect -75 -668 -74 -664
rect -72 -662 -70 -658
rect -66 -662 -64 -658
rect -72 -668 -64 -662
rect -62 -664 -57 -658
rect -62 -668 -61 -664
rect -96 -678 -95 -674
rect -885 -726 -880 -710
rect -881 -730 -880 -726
rect -878 -714 -877 -710
rect -878 -730 -873 -714
rect -861 -726 -856 -710
rect -857 -730 -856 -726
rect -854 -714 -853 -710
rect -854 -730 -849 -714
rect -835 -720 -830 -714
rect -831 -724 -830 -720
rect -828 -718 -827 -714
rect -828 -724 -823 -718
rect -817 -726 -812 -710
rect -813 -730 -812 -726
rect -810 -730 -803 -710
rect -801 -714 -800 -710
rect -801 -730 -796 -714
rect -792 -726 -787 -710
rect -788 -730 -787 -726
rect -785 -730 -778 -710
rect -776 -714 -775 -710
rect 252 -666 253 -662
rect -776 -730 -771 -714
rect -767 -720 -762 -714
rect -763 -724 -762 -720
rect -760 -718 -759 -714
rect -760 -724 -755 -718
rect -600 -715 -594 -711
rect -600 -716 -590 -715
rect -570 -715 -567 -711
rect -577 -716 -567 -715
rect -600 -719 -590 -718
rect -596 -723 -590 -719
rect -577 -719 -567 -718
rect -577 -723 -571 -719
rect 71 -695 76 -689
rect -387 -721 -381 -717
rect -387 -722 -377 -721
rect -357 -721 -354 -717
rect -364 -722 -354 -721
rect -668 -736 -667 -732
rect -672 -742 -667 -736
rect -665 -736 -663 -732
rect -659 -736 -658 -732
rect -665 -742 -658 -736
rect -656 -737 -651 -732
rect -656 -741 -655 -737
rect -656 -742 -651 -741
rect -516 -738 -511 -732
rect -512 -742 -511 -738
rect -509 -736 -508 -732
rect -504 -736 -502 -732
rect -509 -742 -502 -736
rect -500 -736 -499 -732
rect -500 -742 -495 -736
rect -387 -725 -377 -724
rect -383 -729 -377 -725
rect -364 -725 -354 -724
rect -364 -729 -358 -725
rect 75 -699 76 -695
rect 78 -693 80 -689
rect 84 -693 86 -689
rect 78 -699 86 -693
rect 88 -695 93 -689
rect 122 -691 127 -675
rect 126 -695 127 -691
rect 129 -695 137 -675
rect 139 -679 140 -675
rect 139 -695 144 -679
rect 153 -681 158 -675
rect 157 -685 158 -681
rect 160 -679 161 -675
rect 160 -685 165 -679
rect 248 -682 253 -666
rect 255 -682 263 -662
rect 265 -678 270 -662
rect 282 -668 287 -662
rect 286 -672 287 -668
rect 289 -666 291 -662
rect 295 -666 297 -662
rect 289 -672 297 -666
rect 299 -668 304 -662
rect 299 -672 300 -668
rect 332 -666 337 -660
rect 336 -670 337 -666
rect 339 -664 341 -660
rect 345 -664 347 -660
rect 339 -670 347 -664
rect 349 -666 354 -660
rect 369 -661 374 -645
rect 373 -665 374 -661
rect 376 -665 384 -645
rect 386 -649 387 -645
rect 386 -665 391 -649
rect 400 -651 405 -645
rect 404 -655 405 -651
rect 407 -649 408 -645
rect 407 -655 412 -649
rect 445 -665 446 -661
rect 349 -670 350 -666
rect 441 -671 446 -665
rect 448 -667 453 -661
rect 448 -671 449 -667
rect 459 -671 464 -665
rect 463 -675 464 -671
rect 466 -669 468 -665
rect 472 -669 474 -665
rect 466 -675 474 -669
rect 476 -671 481 -665
rect 476 -675 477 -671
rect 265 -682 266 -678
rect 493 -681 498 -665
rect 497 -685 498 -681
rect 500 -685 508 -665
rect 510 -669 511 -665
rect 510 -685 515 -669
rect 524 -671 529 -665
rect 528 -675 529 -671
rect 531 -669 532 -665
rect 531 -675 536 -669
rect 807 -656 812 -640
rect 559 -681 564 -675
rect 563 -685 564 -681
rect 566 -679 568 -675
rect 572 -679 574 -675
rect 566 -685 574 -679
rect 576 -681 581 -675
rect 587 -677 592 -671
rect 591 -681 592 -677
rect 594 -675 595 -671
rect 594 -681 599 -675
rect 811 -660 812 -656
rect 814 -644 815 -640
rect 814 -660 819 -644
rect 831 -656 836 -640
rect 835 -660 836 -656
rect 838 -644 839 -640
rect 838 -660 843 -644
rect 857 -650 862 -644
rect 861 -654 862 -650
rect 864 -648 865 -644
rect 864 -654 869 -648
rect 875 -656 880 -640
rect 879 -660 880 -656
rect 882 -660 889 -640
rect 891 -644 892 -640
rect 891 -660 896 -644
rect 900 -656 905 -640
rect 904 -660 905 -656
rect 907 -660 914 -640
rect 916 -644 917 -640
rect 916 -660 921 -644
rect 925 -650 930 -644
rect 929 -654 930 -650
rect 932 -648 933 -644
rect 932 -654 937 -648
rect 957 -647 962 -641
rect 961 -651 962 -647
rect 964 -645 965 -641
rect 964 -651 969 -645
rect 576 -685 577 -681
rect 618 -693 623 -677
rect 88 -699 89 -695
rect 622 -697 623 -693
rect 625 -697 633 -677
rect 635 -681 636 -677
rect 635 -697 640 -681
rect -99 -723 -93 -719
rect -99 -724 -89 -723
rect -69 -723 -66 -719
rect -76 -724 -66 -723
rect -455 -742 -454 -738
rect -459 -748 -454 -742
rect -452 -742 -450 -738
rect -446 -742 -445 -738
rect -452 -748 -445 -742
rect -443 -744 -438 -738
rect -443 -748 -442 -744
rect -303 -744 -298 -738
rect -299 -748 -298 -744
rect -296 -742 -295 -738
rect -291 -742 -289 -738
rect -296 -748 -289 -742
rect -287 -742 -286 -738
rect -99 -727 -89 -726
rect -95 -731 -89 -727
rect -76 -727 -66 -726
rect -76 -731 -70 -727
rect 262 -727 268 -723
rect 262 -728 272 -727
rect 292 -727 295 -723
rect 285 -728 295 -727
rect -287 -748 -282 -742
rect -167 -744 -166 -740
rect -171 -750 -166 -744
rect -164 -744 -162 -740
rect -158 -744 -157 -740
rect -164 -750 -157 -744
rect -155 -746 -150 -740
rect -155 -750 -154 -746
rect -15 -746 -10 -740
rect -11 -750 -10 -746
rect -8 -744 -7 -740
rect -3 -744 -1 -740
rect -8 -750 -1 -744
rect 1 -744 2 -740
rect 262 -731 272 -730
rect 266 -735 272 -731
rect 285 -731 295 -730
rect 285 -735 291 -731
rect 598 -713 604 -709
rect 598 -714 608 -713
rect 469 -718 485 -714
rect 469 -719 489 -718
rect 469 -729 489 -721
rect 598 -718 608 -716
rect 602 -722 608 -718
rect 598 -724 608 -722
rect 598 -727 608 -726
rect 598 -731 604 -727
rect 469 -732 489 -731
rect 473 -736 489 -732
rect 1 -750 6 -744
rect 194 -748 195 -744
rect 190 -754 195 -748
rect 197 -748 199 -744
rect 203 -748 204 -744
rect 197 -754 204 -748
rect 206 -750 211 -744
rect 206 -754 207 -750
rect 346 -750 351 -744
rect 350 -754 351 -750
rect 353 -748 354 -744
rect 358 -748 360 -744
rect 353 -754 360 -748
rect 362 -748 363 -744
rect 803 -748 808 -732
rect 362 -754 367 -748
rect 469 -752 485 -748
rect 807 -752 808 -748
rect 810 -736 811 -732
rect 810 -752 815 -736
rect 469 -753 489 -752
rect 469 -763 489 -755
rect 827 -748 832 -732
rect 831 -752 832 -748
rect 834 -736 835 -732
rect 834 -752 839 -736
rect 853 -742 858 -736
rect 857 -746 858 -742
rect 860 -740 861 -736
rect 860 -746 865 -740
rect 871 -748 876 -732
rect 875 -752 876 -748
rect 878 -752 885 -732
rect 887 -736 888 -732
rect 887 -752 892 -736
rect 896 -748 901 -732
rect 900 -752 901 -748
rect 903 -752 910 -732
rect 912 -736 913 -732
rect 912 -752 917 -736
rect 921 -742 926 -736
rect 925 -746 926 -742
rect 928 -740 929 -736
rect 928 -746 933 -740
rect 956 -739 961 -733
rect 960 -743 961 -739
rect 963 -737 964 -733
rect 963 -743 968 -737
rect 469 -766 489 -765
rect 473 -770 489 -766
rect -888 -813 -883 -797
rect -884 -817 -883 -813
rect -881 -801 -880 -797
rect -881 -817 -876 -801
rect -864 -813 -859 -797
rect -860 -817 -859 -813
rect -857 -801 -856 -797
rect -857 -817 -852 -801
rect -838 -807 -833 -801
rect -834 -811 -833 -807
rect -831 -805 -830 -801
rect -831 -811 -826 -805
rect -820 -813 -815 -797
rect -816 -817 -815 -813
rect -813 -817 -806 -797
rect -804 -801 -803 -797
rect -804 -817 -799 -801
rect -795 -813 -790 -797
rect -791 -817 -790 -813
rect -788 -817 -781 -797
rect -779 -801 -778 -797
rect -779 -817 -774 -801
rect -770 -807 -765 -801
rect -766 -811 -765 -807
rect -763 -805 -762 -801
rect -763 -811 -758 -805
rect 800 -834 805 -818
rect 804 -838 805 -834
rect 807 -822 808 -818
rect 807 -838 812 -822
rect 824 -834 829 -818
rect 828 -838 829 -834
rect 831 -822 832 -818
rect 831 -838 836 -822
rect 850 -828 855 -822
rect 854 -832 855 -828
rect 857 -826 858 -822
rect 857 -832 862 -826
rect 868 -834 873 -818
rect 872 -838 873 -834
rect 875 -838 882 -818
rect 884 -822 885 -818
rect 884 -838 889 -822
rect 893 -834 898 -818
rect 897 -838 898 -834
rect 900 -838 907 -818
rect 909 -822 910 -818
rect 909 -838 914 -822
rect 918 -828 923 -822
rect 922 -832 923 -828
rect 925 -826 926 -822
rect 925 -832 930 -826
rect 957 -825 962 -819
rect 961 -829 962 -825
rect 964 -823 965 -819
rect 964 -829 969 -823
rect -887 -910 -882 -894
rect -883 -914 -882 -910
rect -880 -898 -879 -894
rect -880 -914 -875 -898
rect -863 -910 -858 -894
rect -859 -914 -858 -910
rect -856 -898 -855 -894
rect -856 -914 -851 -898
rect -837 -904 -832 -898
rect -833 -908 -832 -904
rect -830 -902 -829 -898
rect -830 -908 -825 -902
rect -819 -910 -814 -894
rect -815 -914 -814 -910
rect -812 -914 -805 -894
rect -803 -898 -802 -894
rect -803 -914 -798 -898
rect -794 -910 -789 -894
rect -790 -914 -789 -910
rect -787 -914 -780 -894
rect -778 -898 -777 -894
rect -778 -914 -773 -898
rect -769 -904 -764 -898
rect -765 -908 -764 -904
rect -762 -902 -761 -898
rect -762 -908 -757 -902
rect 801 -931 806 -915
rect 805 -935 806 -931
rect 808 -919 809 -915
rect 808 -935 813 -919
rect 825 -931 830 -915
rect 829 -935 830 -931
rect 832 -919 833 -915
rect 832 -935 837 -919
rect 851 -925 856 -919
rect 855 -929 856 -925
rect 858 -923 859 -919
rect 858 -929 863 -923
rect 869 -931 874 -915
rect 873 -935 874 -931
rect 876 -935 883 -915
rect 885 -919 886 -915
rect 885 -935 890 -919
rect 894 -931 899 -915
rect 898 -935 899 -931
rect 901 -935 908 -915
rect 910 -919 911 -915
rect 910 -935 915 -919
rect 919 -925 924 -919
rect 923 -929 924 -925
rect 926 -923 927 -919
rect 926 -929 931 -923
rect 955 -922 960 -916
rect 959 -926 960 -922
rect 962 -920 963 -916
rect 962 -926 967 -920
rect -889 -1000 -884 -984
rect -885 -1004 -884 -1000
rect -882 -988 -881 -984
rect -882 -1004 -877 -988
rect -865 -1000 -860 -984
rect -861 -1004 -860 -1000
rect -858 -988 -857 -984
rect -858 -1004 -853 -988
rect -839 -994 -834 -988
rect -835 -998 -834 -994
rect -832 -992 -831 -988
rect -832 -998 -827 -992
rect -821 -1000 -816 -984
rect -817 -1004 -816 -1000
rect -814 -1004 -807 -984
rect -805 -988 -804 -984
rect -805 -1004 -800 -988
rect -796 -1000 -791 -984
rect -792 -1004 -791 -1000
rect -789 -1004 -782 -984
rect -780 -988 -779 -984
rect -780 -1004 -775 -988
rect -771 -994 -766 -988
rect -767 -998 -766 -994
rect -764 -992 -763 -988
rect -764 -998 -759 -992
rect -890 -1090 -885 -1074
rect -886 -1094 -885 -1090
rect -883 -1078 -882 -1074
rect -883 -1094 -878 -1078
rect -866 -1090 -861 -1074
rect -862 -1094 -861 -1090
rect -859 -1078 -858 -1074
rect -859 -1094 -854 -1078
rect -840 -1084 -835 -1078
rect -836 -1088 -835 -1084
rect -833 -1082 -832 -1078
rect -833 -1088 -828 -1082
rect -822 -1090 -817 -1074
rect -818 -1094 -817 -1090
rect -815 -1094 -808 -1074
rect -806 -1078 -805 -1074
rect -806 -1094 -801 -1078
rect -797 -1090 -792 -1074
rect -793 -1094 -792 -1090
rect -790 -1094 -783 -1074
rect -781 -1078 -780 -1074
rect -781 -1094 -776 -1078
rect -772 -1084 -767 -1078
rect -768 -1088 -767 -1084
rect -765 -1082 -764 -1078
rect -765 -1088 -760 -1082
rect -891 -1182 -886 -1166
rect -887 -1186 -886 -1182
rect -884 -1170 -883 -1166
rect -884 -1186 -879 -1170
rect -867 -1182 -862 -1166
rect -863 -1186 -862 -1182
rect -860 -1170 -859 -1166
rect -860 -1186 -855 -1170
rect -841 -1176 -836 -1170
rect -837 -1180 -836 -1176
rect -834 -1174 -833 -1170
rect -834 -1180 -829 -1174
rect -823 -1182 -818 -1166
rect -819 -1186 -818 -1182
rect -816 -1186 -809 -1166
rect -807 -1170 -806 -1166
rect -807 -1186 -802 -1170
rect -798 -1182 -793 -1166
rect -794 -1186 -793 -1182
rect -791 -1186 -784 -1166
rect -782 -1170 -781 -1166
rect -782 -1186 -777 -1170
rect -773 -1176 -768 -1170
rect -769 -1180 -768 -1176
rect -766 -1174 -765 -1170
rect -766 -1180 -761 -1174
rect -889 -1278 -884 -1262
rect -885 -1282 -884 -1278
rect -882 -1266 -881 -1262
rect -882 -1282 -877 -1266
rect -865 -1278 -860 -1262
rect -861 -1282 -860 -1278
rect -858 -1266 -857 -1262
rect -858 -1282 -853 -1266
rect -839 -1272 -834 -1266
rect -835 -1276 -834 -1272
rect -832 -1270 -831 -1266
rect -832 -1276 -827 -1270
rect -821 -1278 -816 -1262
rect -817 -1282 -816 -1278
rect -814 -1282 -807 -1262
rect -805 -1266 -804 -1262
rect -805 -1282 -800 -1266
rect -796 -1278 -791 -1262
rect -792 -1282 -791 -1278
rect -789 -1282 -782 -1262
rect -780 -1266 -779 -1262
rect -780 -1282 -775 -1266
rect -771 -1272 -766 -1266
rect -767 -1276 -766 -1272
rect -764 -1270 -763 -1266
rect -764 -1276 -759 -1270
<< pdiffusion >>
rect -875 -504 -874 -500
rect -879 -520 -874 -504
rect -872 -520 -866 -500
rect -864 -516 -859 -500
rect -864 -520 -863 -516
rect -851 -504 -850 -500
rect -855 -520 -850 -504
rect -848 -520 -842 -500
rect -840 -516 -835 -500
rect -840 -520 -839 -516
rect -825 -504 -824 -500
rect -829 -520 -824 -504
rect -822 -516 -817 -500
rect -822 -520 -821 -516
rect -807 -504 -806 -500
rect -811 -520 -806 -504
rect -804 -516 -799 -500
rect -804 -520 -803 -516
rect -782 -504 -781 -500
rect -786 -520 -781 -504
rect -779 -516 -774 -500
rect -779 -520 -778 -516
rect -757 -504 -756 -500
rect -761 -520 -756 -504
rect -754 -516 -749 -500
rect -754 -520 -753 -516
rect 813 -525 814 -521
rect -280 -543 -264 -539
rect 809 -541 814 -525
rect 816 -541 822 -521
rect 824 -537 829 -521
rect 824 -541 825 -537
rect 837 -525 838 -521
rect 833 -541 838 -525
rect 840 -541 846 -521
rect 848 -537 853 -521
rect 848 -541 849 -537
rect 863 -525 864 -521
rect 859 -541 864 -525
rect 866 -537 871 -521
rect 866 -541 867 -537
rect 881 -525 882 -521
rect 877 -541 882 -525
rect 884 -537 889 -521
rect 884 -541 885 -537
rect 906 -525 907 -521
rect 902 -541 907 -525
rect 909 -537 914 -521
rect 909 -541 910 -537
rect 931 -525 932 -521
rect 927 -541 932 -525
rect 934 -537 939 -521
rect 934 -541 935 -537
rect 964 -526 965 -522
rect -284 -544 -264 -543
rect -284 -547 -264 -546
rect -284 -551 -268 -547
rect -208 -555 -207 -551
rect -278 -561 -242 -557
rect -282 -562 -242 -561
rect -282 -572 -242 -564
rect -212 -571 -207 -555
rect -205 -567 -197 -551
rect -205 -571 -203 -567
rect -199 -571 -197 -567
rect -195 -555 -194 -551
rect -195 -571 -190 -555
rect -165 -555 -164 -551
rect -282 -575 -242 -574
rect -282 -579 -246 -575
rect -877 -591 -876 -587
rect -881 -607 -876 -591
rect -874 -607 -868 -587
rect -866 -603 -861 -587
rect -866 -607 -865 -603
rect -853 -591 -852 -587
rect -857 -607 -852 -591
rect -850 -607 -844 -587
rect -842 -603 -837 -587
rect -842 -607 -841 -603
rect -827 -591 -826 -587
rect -831 -607 -826 -591
rect -824 -603 -819 -587
rect -824 -607 -823 -603
rect -809 -591 -808 -587
rect -813 -607 -808 -591
rect -806 -603 -801 -587
rect -806 -607 -805 -603
rect -784 -591 -783 -587
rect -788 -607 -783 -591
rect -781 -603 -776 -587
rect -781 -607 -780 -603
rect -759 -591 -758 -587
rect -763 -607 -758 -591
rect -756 -603 -751 -587
rect -756 -607 -755 -603
rect -576 -596 -575 -592
rect -610 -616 -609 -612
rect -614 -632 -609 -616
rect -607 -628 -599 -612
rect -607 -632 -605 -628
rect -601 -632 -599 -628
rect -597 -616 -596 -612
rect -597 -632 -592 -616
rect -580 -632 -575 -596
rect -573 -632 -565 -592
rect -563 -628 -558 -592
rect -536 -596 -535 -592
rect -540 -612 -535 -596
rect -533 -608 -528 -592
rect -533 -612 -532 -608
rect -512 -596 -511 -592
rect -563 -632 -562 -628
rect -516 -632 -511 -596
rect -509 -632 -501 -592
rect -499 -628 -494 -592
rect -363 -602 -362 -598
rect -499 -632 -498 -628
rect -484 -618 -483 -614
rect -488 -634 -483 -618
rect -481 -630 -476 -614
rect -481 -634 -480 -630
rect -463 -618 -462 -614
rect -467 -634 -462 -618
rect -460 -630 -452 -614
rect -460 -634 -458 -630
rect -454 -634 -452 -630
rect -450 -618 -449 -614
rect -450 -634 -445 -618
rect -397 -622 -396 -618
rect -401 -638 -396 -622
rect -394 -634 -386 -618
rect -394 -638 -392 -634
rect -388 -638 -386 -634
rect -384 -622 -383 -618
rect -384 -638 -379 -622
rect -367 -638 -362 -602
rect -360 -638 -352 -598
rect -350 -634 -345 -598
rect -301 -609 -300 -605
rect -326 -627 -321 -611
rect -322 -631 -321 -627
rect -319 -615 -318 -611
rect -319 -631 -314 -615
rect -305 -625 -300 -609
rect -298 -621 -290 -605
rect -298 -625 -296 -621
rect -292 -625 -290 -621
rect -288 -609 -287 -605
rect -288 -625 -283 -609
rect -350 -638 -349 -634
rect -254 -635 -249 -599
rect -250 -639 -249 -635
rect -247 -639 -239 -599
rect -237 -603 -236 -599
rect -237 -639 -232 -603
rect -169 -591 -164 -555
rect -162 -591 -154 -551
rect -152 -587 -147 -551
rect -152 -591 -151 -587
rect -137 -577 -136 -573
rect -141 -593 -136 -577
rect -134 -589 -129 -573
rect 103 -575 119 -571
rect 103 -576 123 -575
rect 103 -579 123 -578
rect 107 -583 123 -579
rect -134 -593 -133 -589
rect -75 -604 -74 -600
rect -109 -624 -108 -620
rect -113 -640 -108 -624
rect -106 -636 -98 -620
rect -106 -640 -104 -636
rect -100 -640 -98 -636
rect -96 -624 -95 -620
rect -96 -640 -91 -624
rect -79 -640 -74 -604
rect -72 -640 -64 -600
rect -62 -636 -57 -600
rect -32 -621 -27 -605
rect -28 -625 -27 -621
rect -25 -609 -24 -605
rect -25 -625 -20 -609
rect -14 -619 -9 -583
rect -10 -623 -9 -619
rect -7 -623 1 -583
rect 3 -587 4 -583
rect 3 -623 8 -587
rect 33 -587 34 -583
rect 29 -603 34 -587
rect 36 -599 44 -583
rect 36 -603 38 -599
rect 42 -603 44 -599
rect 46 -587 47 -583
rect 960 -542 965 -526
rect 967 -538 972 -522
rect 967 -542 968 -538
rect 46 -603 51 -587
rect 81 -593 117 -589
rect 81 -594 121 -593
rect 81 -604 121 -596
rect 81 -607 121 -606
rect 85 -611 121 -607
rect 286 -608 287 -604
rect -62 -640 -61 -636
rect 252 -628 253 -624
rect 75 -635 76 -631
rect -881 -682 -880 -678
rect -885 -698 -880 -682
rect -878 -698 -872 -678
rect -870 -694 -865 -678
rect -870 -698 -869 -694
rect -857 -682 -856 -678
rect -861 -698 -856 -682
rect -854 -698 -848 -678
rect -846 -694 -841 -678
rect -846 -698 -845 -694
rect -831 -682 -830 -678
rect -835 -698 -830 -682
rect -828 -694 -823 -678
rect -828 -698 -827 -694
rect -813 -682 -812 -678
rect -817 -698 -812 -682
rect -810 -694 -805 -678
rect -810 -698 -809 -694
rect -788 -682 -787 -678
rect -792 -698 -787 -682
rect -785 -694 -780 -678
rect -785 -698 -784 -694
rect -763 -682 -762 -678
rect -767 -698 -762 -682
rect -760 -694 -755 -678
rect 71 -671 76 -635
rect 78 -671 86 -631
rect 88 -667 93 -631
rect 126 -641 127 -637
rect 122 -657 127 -641
rect 129 -653 137 -637
rect 129 -657 131 -653
rect 135 -657 137 -653
rect 139 -641 140 -637
rect 139 -657 144 -641
rect 157 -647 158 -643
rect 88 -671 89 -667
rect -760 -698 -759 -694
rect 153 -663 158 -647
rect 160 -659 165 -643
rect 248 -644 253 -628
rect 255 -640 263 -624
rect 255 -644 257 -640
rect 261 -644 263 -640
rect 265 -628 266 -624
rect 265 -644 270 -628
rect 282 -644 287 -608
rect 289 -644 297 -604
rect 299 -640 304 -604
rect 299 -644 300 -640
rect 336 -606 337 -602
rect 332 -642 337 -606
rect 339 -642 347 -602
rect 349 -638 354 -602
rect 373 -611 374 -607
rect 369 -627 374 -611
rect 376 -623 384 -607
rect 376 -627 378 -623
rect 382 -627 384 -623
rect 386 -611 387 -607
rect 386 -627 391 -611
rect 404 -617 405 -613
rect 349 -642 350 -638
rect 160 -663 161 -659
rect 400 -633 405 -617
rect 407 -629 412 -613
rect 407 -633 408 -629
rect 441 -645 446 -629
rect -672 -715 -667 -699
rect -668 -719 -667 -715
rect -665 -713 -658 -699
rect -665 -717 -663 -713
rect -659 -717 -658 -713
rect -665 -719 -658 -717
rect -656 -703 -655 -699
rect -656 -719 -651 -703
rect -512 -703 -511 -699
rect -627 -715 -612 -710
rect -632 -716 -612 -715
rect -555 -715 -540 -710
rect -555 -716 -535 -715
rect -632 -719 -612 -718
rect -632 -723 -616 -719
rect -555 -719 -535 -718
rect -516 -719 -511 -703
rect -509 -713 -502 -699
rect -509 -717 -508 -713
rect -504 -717 -502 -713
rect -509 -719 -502 -717
rect -500 -715 -495 -699
rect -500 -719 -499 -715
rect -551 -723 -535 -719
rect -459 -721 -454 -705
rect -455 -725 -454 -721
rect -452 -719 -445 -705
rect -452 -723 -450 -719
rect -446 -723 -445 -719
rect -452 -725 -445 -723
rect -443 -709 -442 -705
rect -443 -725 -438 -709
rect -299 -709 -298 -705
rect -414 -721 -399 -716
rect -419 -722 -399 -721
rect -342 -721 -327 -716
rect -342 -722 -322 -721
rect -419 -725 -399 -724
rect -419 -729 -403 -725
rect -342 -725 -322 -724
rect -303 -725 -298 -709
rect -296 -719 -289 -705
rect -296 -723 -295 -719
rect -291 -723 -289 -719
rect -296 -725 -289 -723
rect -287 -721 -282 -705
rect 445 -649 446 -645
rect 448 -633 449 -629
rect 448 -649 453 -633
rect 459 -643 464 -607
rect 463 -647 464 -643
rect 466 -647 474 -607
rect 476 -611 477 -607
rect 476 -647 481 -611
rect 811 -612 812 -608
rect 563 -621 564 -617
rect 497 -631 498 -627
rect 493 -647 498 -631
rect 500 -643 508 -627
rect 500 -647 502 -643
rect 506 -647 508 -643
rect 510 -631 511 -627
rect 510 -647 515 -631
rect 528 -637 529 -633
rect 524 -653 529 -637
rect 531 -649 536 -633
rect 531 -653 532 -649
rect 559 -657 564 -621
rect 566 -657 574 -617
rect 576 -653 581 -617
rect 807 -628 812 -612
rect 814 -628 820 -608
rect 822 -624 827 -608
rect 822 -628 823 -624
rect 835 -612 836 -608
rect 831 -628 836 -612
rect 838 -628 844 -608
rect 846 -624 851 -608
rect 846 -628 847 -624
rect 861 -612 862 -608
rect 857 -628 862 -612
rect 864 -624 869 -608
rect 864 -628 865 -624
rect 879 -612 880 -608
rect 875 -628 880 -612
rect 882 -624 887 -608
rect 882 -628 883 -624
rect 904 -612 905 -608
rect 900 -628 905 -612
rect 907 -624 912 -608
rect 907 -628 908 -624
rect 929 -612 930 -608
rect 925 -628 930 -612
rect 932 -624 937 -608
rect 932 -628 933 -624
rect 961 -613 962 -609
rect 576 -657 577 -653
rect 591 -643 592 -639
rect 587 -659 592 -643
rect 594 -655 599 -639
rect 594 -659 595 -655
rect 622 -643 623 -639
rect 618 -659 623 -643
rect 625 -655 633 -639
rect 625 -659 627 -655
rect 631 -659 633 -655
rect 635 -643 636 -639
rect 635 -659 640 -643
rect 957 -629 962 -613
rect 964 -625 969 -609
rect 964 -629 965 -625
rect -287 -725 -286 -721
rect -171 -723 -166 -707
rect -338 -729 -322 -725
rect -167 -727 -166 -723
rect -164 -721 -157 -707
rect -164 -725 -162 -721
rect -158 -725 -157 -721
rect -164 -727 -157 -725
rect -155 -711 -154 -707
rect -155 -727 -150 -711
rect -11 -711 -10 -707
rect -126 -723 -111 -718
rect -131 -724 -111 -723
rect -54 -723 -39 -718
rect -54 -724 -34 -723
rect -131 -727 -111 -726
rect -131 -731 -115 -727
rect -54 -727 -34 -726
rect -15 -727 -10 -711
rect -8 -721 -1 -707
rect -8 -725 -7 -721
rect -3 -725 -1 -721
rect -8 -727 -1 -725
rect 1 -723 6 -707
rect 807 -704 808 -700
rect 1 -727 2 -723
rect 190 -727 195 -711
rect -50 -731 -34 -727
rect 194 -731 195 -727
rect 197 -725 204 -711
rect 197 -729 199 -725
rect 203 -729 204 -725
rect 197 -731 204 -729
rect 206 -715 207 -711
rect 206 -731 211 -715
rect 350 -715 351 -711
rect 235 -727 250 -722
rect 230 -728 250 -727
rect 307 -727 322 -722
rect 307 -728 327 -727
rect 230 -731 250 -730
rect 230 -735 246 -731
rect 307 -731 327 -730
rect 346 -731 351 -715
rect 353 -725 360 -711
rect 353 -729 354 -725
rect 358 -729 360 -725
rect 353 -731 360 -729
rect 362 -727 367 -711
rect 544 -713 580 -709
rect 540 -714 580 -713
rect 435 -718 451 -714
rect 431 -719 451 -718
rect 362 -731 363 -727
rect 431 -723 451 -721
rect 431 -727 447 -723
rect 431 -729 451 -727
rect 540 -724 580 -716
rect 803 -720 808 -704
rect 810 -720 816 -700
rect 818 -716 823 -700
rect 818 -720 819 -716
rect 831 -704 832 -700
rect 827 -720 832 -704
rect 834 -720 840 -700
rect 842 -716 847 -700
rect 842 -720 843 -716
rect 857 -704 858 -700
rect 853 -720 858 -704
rect 860 -716 865 -700
rect 860 -720 861 -716
rect 875 -704 876 -700
rect 871 -720 876 -704
rect 878 -716 883 -700
rect 878 -720 879 -716
rect 900 -704 901 -700
rect 896 -720 901 -704
rect 903 -716 908 -700
rect 903 -720 904 -716
rect 925 -704 926 -700
rect 921 -720 926 -704
rect 928 -716 933 -700
rect 928 -720 929 -716
rect 960 -705 961 -701
rect 540 -727 580 -726
rect 540 -731 576 -727
rect 311 -735 327 -731
rect 431 -732 451 -731
rect 435 -736 451 -732
rect 435 -752 451 -748
rect 431 -753 451 -752
rect 431 -757 451 -755
rect 431 -761 447 -757
rect 431 -763 451 -761
rect 956 -721 961 -705
rect 963 -717 968 -701
rect 963 -721 964 -717
rect -884 -769 -883 -765
rect -888 -785 -883 -769
rect -881 -785 -875 -765
rect -873 -781 -868 -765
rect -873 -785 -872 -781
rect -860 -769 -859 -765
rect -864 -785 -859 -769
rect -857 -785 -851 -765
rect -849 -781 -844 -765
rect -849 -785 -848 -781
rect -834 -769 -833 -765
rect -838 -785 -833 -769
rect -831 -781 -826 -765
rect -831 -785 -830 -781
rect -816 -769 -815 -765
rect -820 -785 -815 -769
rect -813 -781 -808 -765
rect -813 -785 -812 -781
rect -791 -769 -790 -765
rect -795 -785 -790 -769
rect -788 -781 -783 -765
rect -788 -785 -787 -781
rect -766 -769 -765 -765
rect -770 -785 -765 -769
rect -763 -781 -758 -765
rect 431 -766 451 -765
rect 435 -770 451 -766
rect -763 -785 -762 -781
rect 804 -790 805 -786
rect 800 -806 805 -790
rect 807 -806 813 -786
rect 815 -802 820 -786
rect 815 -806 816 -802
rect 828 -790 829 -786
rect 824 -806 829 -790
rect 831 -806 837 -786
rect 839 -802 844 -786
rect 839 -806 840 -802
rect 854 -790 855 -786
rect 850 -806 855 -790
rect 857 -802 862 -786
rect 857 -806 858 -802
rect 872 -790 873 -786
rect 868 -806 873 -790
rect 875 -802 880 -786
rect 875 -806 876 -802
rect 897 -790 898 -786
rect 893 -806 898 -790
rect 900 -802 905 -786
rect 900 -806 901 -802
rect 922 -790 923 -786
rect 918 -806 923 -790
rect 925 -802 930 -786
rect 925 -806 926 -802
rect 961 -791 962 -787
rect 957 -807 962 -791
rect 964 -803 969 -787
rect 964 -807 965 -803
rect -883 -866 -882 -862
rect -887 -882 -882 -866
rect -880 -882 -874 -862
rect -872 -878 -867 -862
rect -872 -882 -871 -878
rect -859 -866 -858 -862
rect -863 -882 -858 -866
rect -856 -882 -850 -862
rect -848 -878 -843 -862
rect -848 -882 -847 -878
rect -833 -866 -832 -862
rect -837 -882 -832 -866
rect -830 -878 -825 -862
rect -830 -882 -829 -878
rect -815 -866 -814 -862
rect -819 -882 -814 -866
rect -812 -878 -807 -862
rect -812 -882 -811 -878
rect -790 -866 -789 -862
rect -794 -882 -789 -866
rect -787 -878 -782 -862
rect -787 -882 -786 -878
rect -765 -866 -764 -862
rect -769 -882 -764 -866
rect -762 -878 -757 -862
rect -762 -882 -761 -878
rect 805 -887 806 -883
rect 801 -903 806 -887
rect 808 -903 814 -883
rect 816 -899 821 -883
rect 816 -903 817 -899
rect 829 -887 830 -883
rect 825 -903 830 -887
rect 832 -903 838 -883
rect 840 -899 845 -883
rect 840 -903 841 -899
rect 855 -887 856 -883
rect 851 -903 856 -887
rect 858 -899 863 -883
rect 858 -903 859 -899
rect 873 -887 874 -883
rect 869 -903 874 -887
rect 876 -899 881 -883
rect 876 -903 877 -899
rect 898 -887 899 -883
rect 894 -903 899 -887
rect 901 -899 906 -883
rect 901 -903 902 -899
rect 923 -887 924 -883
rect 919 -903 924 -887
rect 926 -899 931 -883
rect 926 -903 927 -899
rect 959 -888 960 -884
rect 955 -904 960 -888
rect 962 -900 967 -884
rect 962 -904 963 -900
rect -885 -956 -884 -952
rect -889 -972 -884 -956
rect -882 -972 -876 -952
rect -874 -968 -869 -952
rect -874 -972 -873 -968
rect -861 -956 -860 -952
rect -865 -972 -860 -956
rect -858 -972 -852 -952
rect -850 -968 -845 -952
rect -850 -972 -849 -968
rect -835 -956 -834 -952
rect -839 -972 -834 -956
rect -832 -968 -827 -952
rect -832 -972 -831 -968
rect -817 -956 -816 -952
rect -821 -972 -816 -956
rect -814 -968 -809 -952
rect -814 -972 -813 -968
rect -792 -956 -791 -952
rect -796 -972 -791 -956
rect -789 -968 -784 -952
rect -789 -972 -788 -968
rect -767 -956 -766 -952
rect -771 -972 -766 -956
rect -764 -968 -759 -952
rect -764 -972 -763 -968
rect -886 -1046 -885 -1042
rect -890 -1062 -885 -1046
rect -883 -1062 -877 -1042
rect -875 -1058 -870 -1042
rect -875 -1062 -874 -1058
rect -862 -1046 -861 -1042
rect -866 -1062 -861 -1046
rect -859 -1062 -853 -1042
rect -851 -1058 -846 -1042
rect -851 -1062 -850 -1058
rect -836 -1046 -835 -1042
rect -840 -1062 -835 -1046
rect -833 -1058 -828 -1042
rect -833 -1062 -832 -1058
rect -818 -1046 -817 -1042
rect -822 -1062 -817 -1046
rect -815 -1058 -810 -1042
rect -815 -1062 -814 -1058
rect -793 -1046 -792 -1042
rect -797 -1062 -792 -1046
rect -790 -1058 -785 -1042
rect -790 -1062 -789 -1058
rect -768 -1046 -767 -1042
rect -772 -1062 -767 -1046
rect -765 -1058 -760 -1042
rect -765 -1062 -764 -1058
rect -887 -1138 -886 -1134
rect -891 -1154 -886 -1138
rect -884 -1154 -878 -1134
rect -876 -1150 -871 -1134
rect -876 -1154 -875 -1150
rect -863 -1138 -862 -1134
rect -867 -1154 -862 -1138
rect -860 -1154 -854 -1134
rect -852 -1150 -847 -1134
rect -852 -1154 -851 -1150
rect -837 -1138 -836 -1134
rect -841 -1154 -836 -1138
rect -834 -1150 -829 -1134
rect -834 -1154 -833 -1150
rect -819 -1138 -818 -1134
rect -823 -1154 -818 -1138
rect -816 -1150 -811 -1134
rect -816 -1154 -815 -1150
rect -794 -1138 -793 -1134
rect -798 -1154 -793 -1138
rect -791 -1150 -786 -1134
rect -791 -1154 -790 -1150
rect -769 -1138 -768 -1134
rect -773 -1154 -768 -1138
rect -766 -1150 -761 -1134
rect -766 -1154 -765 -1150
rect -885 -1234 -884 -1230
rect -889 -1250 -884 -1234
rect -882 -1250 -876 -1230
rect -874 -1246 -869 -1230
rect -874 -1250 -873 -1246
rect -861 -1234 -860 -1230
rect -865 -1250 -860 -1234
rect -858 -1250 -852 -1230
rect -850 -1246 -845 -1230
rect -850 -1250 -849 -1246
rect -835 -1234 -834 -1230
rect -839 -1250 -834 -1234
rect -832 -1246 -827 -1230
rect -832 -1250 -831 -1246
rect -817 -1234 -816 -1230
rect -821 -1250 -816 -1234
rect -814 -1246 -809 -1230
rect -814 -1250 -813 -1246
rect -792 -1234 -791 -1230
rect -796 -1250 -791 -1234
rect -789 -1246 -784 -1230
rect -789 -1250 -788 -1246
rect -767 -1234 -766 -1230
rect -771 -1250 -766 -1234
rect -764 -1246 -759 -1230
rect -764 -1250 -763 -1246
<< ndcontact >>
rect -879 -552 -875 -548
rect -871 -536 -867 -532
rect -855 -552 -851 -548
rect -847 -536 -843 -532
rect -829 -546 -825 -542
rect -821 -540 -817 -536
rect -811 -552 -807 -548
rect -794 -536 -790 -532
rect -786 -552 -782 -548
rect -769 -536 -765 -532
rect -761 -546 -757 -542
rect -753 -540 -749 -536
rect -300 -543 -296 -539
rect -306 -551 -302 -547
rect -310 -561 -306 -557
rect -304 -570 -300 -566
rect -310 -579 -306 -575
rect -881 -639 -877 -635
rect -873 -623 -869 -619
rect -857 -639 -853 -635
rect -849 -623 -845 -619
rect -831 -633 -827 -629
rect -823 -627 -819 -623
rect -813 -639 -809 -635
rect -796 -623 -792 -619
rect -788 -639 -784 -635
rect -771 -623 -767 -619
rect -763 -633 -759 -629
rect -755 -627 -751 -623
rect -540 -634 -536 -630
rect -532 -628 -528 -624
rect -614 -654 -610 -650
rect -580 -660 -576 -656
rect -571 -654 -567 -650
rect -562 -660 -558 -656
rect -516 -660 -512 -656
rect -507 -654 -503 -650
rect -488 -656 -484 -652
rect -480 -650 -476 -646
rect -498 -660 -494 -656
rect -596 -670 -592 -666
rect -467 -672 -463 -668
rect -449 -656 -445 -652
rect -212 -609 -208 -605
rect -194 -593 -190 -589
rect 135 -575 139 -571
rect 809 -573 813 -569
rect 817 -557 821 -553
rect 141 -583 145 -579
rect 833 -573 837 -569
rect 841 -557 845 -553
rect -169 -619 -165 -615
rect -160 -613 -156 -609
rect -141 -615 -137 -611
rect -133 -609 -129 -605
rect -151 -619 -147 -615
rect -326 -647 -322 -643
rect -318 -653 -314 -649
rect -305 -647 -301 -643
rect -401 -660 -397 -656
rect -367 -666 -363 -662
rect -358 -660 -354 -656
rect -349 -666 -345 -662
rect 859 -567 863 -563
rect 867 -561 871 -557
rect 877 -573 881 -569
rect 894 -557 898 -553
rect 902 -573 906 -569
rect 919 -557 923 -553
rect 927 -567 931 -563
rect 935 -561 939 -557
rect 960 -564 964 -560
rect 968 -558 972 -554
rect 145 -593 149 -589
rect 139 -602 143 -598
rect 145 -611 149 -607
rect -287 -663 -283 -659
rect -254 -667 -250 -663
rect -245 -661 -241 -657
rect -32 -641 -28 -637
rect 29 -625 33 -621
rect 47 -641 51 -637
rect -24 -647 -20 -643
rect -14 -651 -10 -647
rect -5 -645 -1 -641
rect 4 -651 8 -647
rect -236 -667 -232 -663
rect -113 -662 -109 -658
rect -383 -676 -379 -672
rect -79 -668 -75 -664
rect -70 -662 -66 -658
rect -61 -668 -57 -664
rect -95 -678 -91 -674
rect -885 -730 -881 -726
rect -877 -714 -873 -710
rect -861 -730 -857 -726
rect -853 -714 -849 -710
rect -835 -724 -831 -720
rect -827 -718 -823 -714
rect -817 -730 -813 -726
rect -800 -714 -796 -710
rect -792 -730 -788 -726
rect -775 -714 -771 -710
rect 248 -666 252 -662
rect -767 -724 -763 -720
rect -759 -718 -755 -714
rect -594 -715 -590 -711
rect -577 -715 -570 -711
rect -600 -723 -596 -719
rect -571 -723 -567 -719
rect -381 -721 -377 -717
rect -364 -721 -357 -717
rect -672 -736 -668 -732
rect -663 -736 -659 -732
rect -655 -741 -651 -737
rect -516 -742 -512 -738
rect -508 -736 -504 -732
rect -499 -736 -495 -732
rect -387 -729 -383 -725
rect -358 -729 -354 -725
rect 71 -699 75 -695
rect 80 -693 84 -689
rect 122 -695 126 -691
rect 140 -679 144 -675
rect 153 -685 157 -681
rect 161 -679 165 -675
rect 282 -672 286 -668
rect 291 -666 295 -662
rect 300 -672 304 -668
rect 332 -670 336 -666
rect 341 -664 345 -660
rect 369 -665 373 -661
rect 387 -649 391 -645
rect 400 -655 404 -651
rect 408 -649 412 -645
rect 441 -665 445 -661
rect 350 -670 354 -666
rect 449 -671 453 -667
rect 459 -675 463 -671
rect 468 -669 472 -665
rect 477 -675 481 -671
rect 266 -682 270 -678
rect 493 -685 497 -681
rect 511 -669 515 -665
rect 524 -675 528 -671
rect 532 -669 536 -665
rect 559 -685 563 -681
rect 568 -679 572 -675
rect 587 -681 591 -677
rect 595 -675 599 -671
rect 807 -660 811 -656
rect 815 -644 819 -640
rect 831 -660 835 -656
rect 839 -644 843 -640
rect 857 -654 861 -650
rect 865 -648 869 -644
rect 875 -660 879 -656
rect 892 -644 896 -640
rect 900 -660 904 -656
rect 917 -644 921 -640
rect 925 -654 929 -650
rect 933 -648 937 -644
rect 957 -651 961 -647
rect 965 -645 969 -641
rect 577 -685 581 -681
rect 89 -699 93 -695
rect 618 -697 622 -693
rect 636 -681 640 -677
rect -93 -723 -89 -719
rect -76 -723 -69 -719
rect -459 -742 -455 -738
rect -450 -742 -446 -738
rect -442 -748 -438 -744
rect -303 -748 -299 -744
rect -295 -742 -291 -738
rect -286 -742 -282 -738
rect -99 -731 -95 -727
rect -70 -731 -66 -727
rect 268 -727 272 -723
rect 285 -727 292 -723
rect -171 -744 -167 -740
rect -162 -744 -158 -740
rect -154 -750 -150 -746
rect -15 -750 -11 -746
rect -7 -744 -3 -740
rect 2 -744 6 -740
rect 262 -735 266 -731
rect 291 -735 295 -731
rect 604 -713 608 -709
rect 485 -718 489 -714
rect 598 -722 602 -718
rect 604 -731 608 -727
rect 469 -736 473 -732
rect 190 -748 194 -744
rect 199 -748 203 -744
rect 207 -754 211 -750
rect 346 -754 350 -750
rect 354 -748 358 -744
rect 363 -748 367 -744
rect 485 -752 489 -748
rect 803 -752 807 -748
rect 811 -736 815 -732
rect 827 -752 831 -748
rect 835 -736 839 -732
rect 853 -746 857 -742
rect 861 -740 865 -736
rect 871 -752 875 -748
rect 888 -736 892 -732
rect 896 -752 900 -748
rect 913 -736 917 -732
rect 921 -746 925 -742
rect 929 -740 933 -736
rect 956 -743 960 -739
rect 964 -737 968 -733
rect 469 -770 473 -766
rect -888 -817 -884 -813
rect -880 -801 -876 -797
rect -864 -817 -860 -813
rect -856 -801 -852 -797
rect -838 -811 -834 -807
rect -830 -805 -826 -801
rect -820 -817 -816 -813
rect -803 -801 -799 -797
rect -795 -817 -791 -813
rect -778 -801 -774 -797
rect -770 -811 -766 -807
rect -762 -805 -758 -801
rect 800 -838 804 -834
rect 808 -822 812 -818
rect 824 -838 828 -834
rect 832 -822 836 -818
rect 850 -832 854 -828
rect 858 -826 862 -822
rect 868 -838 872 -834
rect 885 -822 889 -818
rect 893 -838 897 -834
rect 910 -822 914 -818
rect 918 -832 922 -828
rect 926 -826 930 -822
rect 957 -829 961 -825
rect 965 -823 969 -819
rect -887 -914 -883 -910
rect -879 -898 -875 -894
rect -863 -914 -859 -910
rect -855 -898 -851 -894
rect -837 -908 -833 -904
rect -829 -902 -825 -898
rect -819 -914 -815 -910
rect -802 -898 -798 -894
rect -794 -914 -790 -910
rect -777 -898 -773 -894
rect -769 -908 -765 -904
rect -761 -902 -757 -898
rect 801 -935 805 -931
rect 809 -919 813 -915
rect 825 -935 829 -931
rect 833 -919 837 -915
rect 851 -929 855 -925
rect 859 -923 863 -919
rect 869 -935 873 -931
rect 886 -919 890 -915
rect 894 -935 898 -931
rect 911 -919 915 -915
rect 919 -929 923 -925
rect 927 -923 931 -919
rect 955 -926 959 -922
rect 963 -920 967 -916
rect -889 -1004 -885 -1000
rect -881 -988 -877 -984
rect -865 -1004 -861 -1000
rect -857 -988 -853 -984
rect -839 -998 -835 -994
rect -831 -992 -827 -988
rect -821 -1004 -817 -1000
rect -804 -988 -800 -984
rect -796 -1004 -792 -1000
rect -779 -988 -775 -984
rect -771 -998 -767 -994
rect -763 -992 -759 -988
rect -890 -1094 -886 -1090
rect -882 -1078 -878 -1074
rect -866 -1094 -862 -1090
rect -858 -1078 -854 -1074
rect -840 -1088 -836 -1084
rect -832 -1082 -828 -1078
rect -822 -1094 -818 -1090
rect -805 -1078 -801 -1074
rect -797 -1094 -793 -1090
rect -780 -1078 -776 -1074
rect -772 -1088 -768 -1084
rect -764 -1082 -760 -1078
rect -891 -1186 -887 -1182
rect -883 -1170 -879 -1166
rect -867 -1186 -863 -1182
rect -859 -1170 -855 -1166
rect -841 -1180 -837 -1176
rect -833 -1174 -829 -1170
rect -823 -1186 -819 -1182
rect -806 -1170 -802 -1166
rect -798 -1186 -794 -1182
rect -781 -1170 -777 -1166
rect -773 -1180 -769 -1176
rect -765 -1174 -761 -1170
rect -889 -1282 -885 -1278
rect -881 -1266 -877 -1262
rect -865 -1282 -861 -1278
rect -857 -1266 -853 -1262
rect -839 -1276 -835 -1272
rect -831 -1270 -827 -1266
rect -821 -1282 -817 -1278
rect -804 -1266 -800 -1262
rect -796 -1282 -792 -1278
rect -779 -1266 -775 -1262
rect -771 -1276 -767 -1272
rect -763 -1270 -759 -1266
<< pdcontact >>
rect -879 -504 -875 -500
rect -863 -520 -859 -516
rect -855 -504 -851 -500
rect -839 -520 -835 -516
rect -829 -504 -825 -500
rect -821 -520 -817 -516
rect -811 -504 -807 -500
rect -803 -520 -799 -516
rect -786 -504 -782 -500
rect -778 -520 -774 -516
rect -761 -504 -757 -500
rect -753 -520 -749 -516
rect 809 -525 813 -521
rect -284 -543 -280 -539
rect 825 -541 829 -537
rect 833 -525 837 -521
rect 849 -541 853 -537
rect 859 -525 863 -521
rect 867 -541 871 -537
rect 877 -525 881 -521
rect 885 -541 889 -537
rect 902 -525 906 -521
rect 910 -541 914 -537
rect 927 -525 931 -521
rect 935 -541 939 -537
rect 960 -526 964 -522
rect -268 -551 -264 -547
rect -212 -555 -208 -551
rect -282 -561 -278 -557
rect -203 -571 -199 -567
rect -194 -555 -190 -551
rect -169 -555 -165 -551
rect -246 -579 -242 -575
rect -881 -591 -877 -587
rect -865 -607 -861 -603
rect -857 -591 -853 -587
rect -841 -607 -837 -603
rect -831 -591 -827 -587
rect -823 -607 -819 -603
rect -813 -591 -809 -587
rect -805 -607 -801 -603
rect -788 -591 -784 -587
rect -780 -607 -776 -603
rect -763 -591 -759 -587
rect -755 -607 -751 -603
rect -580 -596 -576 -592
rect -614 -616 -610 -612
rect -605 -632 -601 -628
rect -596 -616 -592 -612
rect -540 -596 -536 -592
rect -532 -612 -528 -608
rect -516 -596 -512 -592
rect -562 -632 -558 -628
rect -367 -602 -363 -598
rect -498 -632 -494 -628
rect -488 -618 -484 -614
rect -480 -634 -476 -630
rect -467 -618 -463 -614
rect -458 -634 -454 -630
rect -449 -618 -445 -614
rect -401 -622 -397 -618
rect -392 -638 -388 -634
rect -383 -622 -379 -618
rect -305 -609 -301 -605
rect -326 -631 -322 -627
rect -318 -615 -314 -611
rect -296 -625 -292 -621
rect -287 -609 -283 -605
rect -349 -638 -345 -634
rect -254 -639 -250 -635
rect -236 -603 -232 -599
rect -151 -591 -147 -587
rect -141 -577 -137 -573
rect 119 -575 123 -571
rect 103 -583 107 -579
rect -133 -593 -129 -589
rect -79 -604 -75 -600
rect -113 -624 -109 -620
rect -104 -640 -100 -636
rect -95 -624 -91 -620
rect -32 -625 -28 -621
rect -24 -609 -20 -605
rect -14 -623 -10 -619
rect 4 -587 8 -583
rect 29 -587 33 -583
rect 38 -603 42 -599
rect 47 -587 51 -583
rect 968 -542 972 -538
rect 117 -593 121 -589
rect 81 -611 85 -607
rect 282 -608 286 -604
rect -61 -640 -57 -636
rect 248 -628 252 -624
rect 71 -635 75 -631
rect -885 -682 -881 -678
rect -869 -698 -865 -694
rect -861 -682 -857 -678
rect -845 -698 -841 -694
rect -835 -682 -831 -678
rect -827 -698 -823 -694
rect -817 -682 -813 -678
rect -809 -698 -805 -694
rect -792 -682 -788 -678
rect -784 -698 -780 -694
rect -767 -682 -763 -678
rect 122 -641 126 -637
rect 131 -657 135 -653
rect 140 -641 144 -637
rect 153 -647 157 -643
rect 89 -671 93 -667
rect -759 -698 -755 -694
rect 257 -644 261 -640
rect 266 -628 270 -624
rect 300 -644 304 -640
rect 332 -606 336 -602
rect 369 -611 373 -607
rect 378 -627 382 -623
rect 387 -611 391 -607
rect 400 -617 404 -613
rect 350 -642 354 -638
rect 161 -663 165 -659
rect 408 -633 412 -629
rect -672 -719 -668 -715
rect -663 -717 -659 -713
rect -655 -703 -651 -699
rect -516 -703 -512 -699
rect -616 -723 -612 -719
rect -508 -717 -504 -713
rect -499 -719 -495 -715
rect -555 -723 -551 -719
rect -459 -725 -455 -721
rect -450 -723 -446 -719
rect -442 -709 -438 -705
rect -303 -709 -299 -705
rect -403 -729 -399 -725
rect -295 -723 -291 -719
rect 441 -649 445 -645
rect 449 -633 453 -629
rect 459 -647 463 -643
rect 477 -611 481 -607
rect 807 -612 811 -608
rect 559 -621 563 -617
rect 493 -631 497 -627
rect 502 -647 506 -643
rect 511 -631 515 -627
rect 524 -637 528 -633
rect 532 -653 536 -649
rect 823 -628 827 -624
rect 831 -612 835 -608
rect 847 -628 851 -624
rect 857 -612 861 -608
rect 865 -628 869 -624
rect 875 -612 879 -608
rect 883 -628 887 -624
rect 900 -612 904 -608
rect 908 -628 912 -624
rect 925 -612 929 -608
rect 933 -628 937 -624
rect 957 -613 961 -609
rect 577 -657 581 -653
rect 587 -643 591 -639
rect 595 -659 599 -655
rect 618 -643 622 -639
rect 627 -659 631 -655
rect 636 -643 640 -639
rect 965 -629 969 -625
rect -286 -725 -282 -721
rect -342 -729 -338 -725
rect -171 -727 -167 -723
rect -162 -725 -158 -721
rect -154 -711 -150 -707
rect -15 -711 -11 -707
rect -115 -731 -111 -727
rect -7 -725 -3 -721
rect 803 -704 807 -700
rect 2 -727 6 -723
rect -54 -731 -50 -727
rect 190 -731 194 -727
rect 199 -729 203 -725
rect 207 -715 211 -711
rect 346 -715 350 -711
rect 246 -735 250 -731
rect 354 -729 358 -725
rect 540 -713 544 -709
rect 431 -718 435 -714
rect 363 -731 367 -727
rect 447 -727 451 -723
rect 819 -720 823 -716
rect 827 -704 831 -700
rect 843 -720 847 -716
rect 853 -704 857 -700
rect 861 -720 865 -716
rect 871 -704 875 -700
rect 879 -720 883 -716
rect 896 -704 900 -700
rect 904 -720 908 -716
rect 921 -704 925 -700
rect 929 -720 933 -716
rect 956 -705 960 -701
rect 576 -731 580 -727
rect 307 -735 311 -731
rect 431 -736 435 -732
rect 431 -752 435 -748
rect 447 -761 451 -757
rect 964 -721 968 -717
rect -888 -769 -884 -765
rect -872 -785 -868 -781
rect -864 -769 -860 -765
rect -848 -785 -844 -781
rect -838 -769 -834 -765
rect -830 -785 -826 -781
rect -820 -769 -816 -765
rect -812 -785 -808 -781
rect -795 -769 -791 -765
rect -787 -785 -783 -781
rect -770 -769 -766 -765
rect 431 -770 435 -766
rect -762 -785 -758 -781
rect 800 -790 804 -786
rect 816 -806 820 -802
rect 824 -790 828 -786
rect 840 -806 844 -802
rect 850 -790 854 -786
rect 858 -806 862 -802
rect 868 -790 872 -786
rect 876 -806 880 -802
rect 893 -790 897 -786
rect 901 -806 905 -802
rect 918 -790 922 -786
rect 926 -806 930 -802
rect 957 -791 961 -787
rect 965 -807 969 -803
rect -887 -866 -883 -862
rect -871 -882 -867 -878
rect -863 -866 -859 -862
rect -847 -882 -843 -878
rect -837 -866 -833 -862
rect -829 -882 -825 -878
rect -819 -866 -815 -862
rect -811 -882 -807 -878
rect -794 -866 -790 -862
rect -786 -882 -782 -878
rect -769 -866 -765 -862
rect -761 -882 -757 -878
rect 801 -887 805 -883
rect 817 -903 821 -899
rect 825 -887 829 -883
rect 841 -903 845 -899
rect 851 -887 855 -883
rect 859 -903 863 -899
rect 869 -887 873 -883
rect 877 -903 881 -899
rect 894 -887 898 -883
rect 902 -903 906 -899
rect 919 -887 923 -883
rect 927 -903 931 -899
rect 955 -888 959 -884
rect 963 -904 967 -900
rect -889 -956 -885 -952
rect -873 -972 -869 -968
rect -865 -956 -861 -952
rect -849 -972 -845 -968
rect -839 -956 -835 -952
rect -831 -972 -827 -968
rect -821 -956 -817 -952
rect -813 -972 -809 -968
rect -796 -956 -792 -952
rect -788 -972 -784 -968
rect -771 -956 -767 -952
rect -763 -972 -759 -968
rect -890 -1046 -886 -1042
rect -874 -1062 -870 -1058
rect -866 -1046 -862 -1042
rect -850 -1062 -846 -1058
rect -840 -1046 -836 -1042
rect -832 -1062 -828 -1058
rect -822 -1046 -818 -1042
rect -814 -1062 -810 -1058
rect -797 -1046 -793 -1042
rect -789 -1062 -785 -1058
rect -772 -1046 -768 -1042
rect -764 -1062 -760 -1058
rect -891 -1138 -887 -1134
rect -875 -1154 -871 -1150
rect -867 -1138 -863 -1134
rect -851 -1154 -847 -1150
rect -841 -1138 -837 -1134
rect -833 -1154 -829 -1150
rect -823 -1138 -819 -1134
rect -815 -1154 -811 -1150
rect -798 -1138 -794 -1134
rect -790 -1154 -786 -1150
rect -773 -1138 -769 -1134
rect -765 -1154 -761 -1150
rect -889 -1234 -885 -1230
rect -873 -1250 -869 -1246
rect -865 -1234 -861 -1230
rect -849 -1250 -845 -1246
rect -839 -1234 -835 -1230
rect -831 -1250 -827 -1246
rect -821 -1234 -817 -1230
rect -813 -1250 -809 -1246
rect -796 -1234 -792 -1230
rect -788 -1250 -784 -1246
rect -771 -1234 -767 -1230
rect -763 -1250 -759 -1246
<< polysilicon >>
rect -874 -500 -872 -496
rect -866 -500 -864 -496
rect -850 -500 -848 -496
rect -842 -500 -840 -496
rect -824 -500 -822 -496
rect -806 -500 -804 -497
rect -781 -500 -779 -497
rect -756 -500 -754 -496
rect -874 -532 -872 -520
rect -874 -555 -872 -552
rect -866 -561 -864 -520
rect -850 -532 -848 -520
rect -850 -555 -848 -552
rect -865 -564 -864 -561
rect -842 -564 -840 -520
rect -824 -536 -822 -520
rect -806 -532 -804 -520
rect -797 -532 -795 -528
rect -781 -532 -779 -520
rect -772 -532 -770 -528
rect -824 -550 -822 -546
rect -756 -536 -754 -520
rect 814 -521 816 -517
rect 822 -521 824 -517
rect 838 -521 840 -517
rect 846 -521 848 -517
rect 864 -521 866 -517
rect 882 -521 884 -518
rect 907 -521 909 -518
rect 932 -521 934 -517
rect 965 -522 967 -518
rect -309 -546 -306 -544
rect -296 -546 -284 -544
rect -264 -546 -261 -544
rect -756 -550 -754 -546
rect -207 -551 -205 -547
rect -197 -551 -195 -547
rect -164 -551 -162 -548
rect -154 -551 -152 -548
rect -806 -557 -804 -552
rect -797 -566 -795 -552
rect -781 -557 -779 -552
rect -772 -566 -770 -552
rect -313 -564 -310 -562
rect -300 -564 -282 -562
rect -242 -564 -239 -562
rect -313 -574 -310 -572
rect -300 -574 -282 -572
rect -242 -574 -239 -572
rect -876 -587 -874 -583
rect -868 -587 -866 -583
rect -852 -587 -850 -583
rect -844 -587 -842 -583
rect -826 -587 -824 -583
rect -808 -587 -806 -584
rect -783 -587 -781 -584
rect -758 -587 -756 -583
rect -575 -592 -573 -589
rect -565 -592 -563 -589
rect -535 -592 -533 -588
rect -207 -589 -205 -571
rect -197 -589 -195 -571
rect -511 -592 -509 -589
rect -501 -592 -499 -589
rect -876 -619 -874 -607
rect -876 -642 -874 -639
rect -868 -648 -866 -607
rect -852 -619 -850 -607
rect -852 -642 -850 -639
rect -867 -651 -866 -648
rect -844 -651 -842 -607
rect -826 -623 -824 -607
rect -808 -619 -806 -607
rect -799 -619 -797 -615
rect -783 -619 -781 -607
rect -774 -619 -772 -615
rect -826 -637 -824 -633
rect -758 -623 -756 -607
rect -609 -612 -607 -608
rect -599 -612 -597 -608
rect -535 -624 -533 -612
rect -758 -637 -756 -633
rect -808 -644 -806 -639
rect -799 -653 -797 -639
rect -783 -644 -781 -639
rect -774 -653 -772 -639
rect -609 -650 -607 -632
rect -599 -650 -597 -632
rect -575 -650 -573 -632
rect -565 -650 -563 -632
rect -362 -598 -360 -595
rect -352 -598 -350 -595
rect -483 -614 -481 -611
rect -462 -614 -460 -610
rect -452 -614 -450 -610
rect -535 -638 -533 -634
rect -511 -650 -509 -632
rect -501 -650 -499 -632
rect -396 -618 -394 -614
rect -386 -618 -384 -614
rect -483 -646 -481 -634
rect -462 -652 -460 -634
rect -452 -652 -450 -634
rect -249 -599 -247 -596
rect -239 -599 -237 -596
rect -300 -605 -298 -601
rect -290 -605 -288 -601
rect -321 -611 -319 -607
rect -483 -659 -481 -656
rect -575 -663 -573 -660
rect -565 -663 -563 -660
rect -511 -663 -509 -660
rect -501 -663 -499 -660
rect -609 -674 -607 -670
rect -599 -674 -597 -670
rect -396 -656 -394 -638
rect -386 -656 -384 -638
rect -362 -656 -360 -638
rect -352 -656 -350 -638
rect -321 -643 -319 -631
rect -300 -643 -298 -625
rect -290 -643 -288 -625
rect 814 -553 816 -541
rect -136 -573 -134 -570
rect -164 -609 -162 -591
rect -154 -609 -152 -591
rect 814 -576 816 -573
rect 100 -578 103 -576
rect 123 -578 135 -576
rect 145 -578 148 -576
rect -9 -583 -7 -580
rect 1 -583 3 -580
rect 34 -583 36 -579
rect 44 -583 46 -579
rect 822 -582 824 -541
rect 838 -553 840 -541
rect 838 -576 840 -573
rect -136 -605 -134 -593
rect -74 -600 -72 -597
rect -64 -600 -62 -597
rect -207 -613 -205 -609
rect -197 -613 -195 -609
rect -136 -618 -134 -615
rect -164 -622 -162 -619
rect -154 -622 -152 -619
rect -108 -620 -106 -616
rect -98 -620 -96 -616
rect -880 -678 -878 -674
rect -872 -678 -870 -674
rect -856 -678 -854 -674
rect -848 -678 -846 -674
rect -830 -678 -828 -674
rect -812 -678 -810 -675
rect -787 -678 -785 -675
rect -762 -678 -760 -674
rect -462 -676 -460 -672
rect -452 -676 -450 -672
rect -321 -657 -319 -653
rect -249 -657 -247 -639
rect -239 -657 -237 -639
rect -27 -605 -25 -602
rect 823 -585 824 -582
rect 846 -585 848 -541
rect 864 -557 866 -541
rect 882 -553 884 -541
rect 891 -553 893 -549
rect 907 -553 909 -541
rect 916 -553 918 -549
rect 864 -571 866 -567
rect 932 -557 934 -541
rect 965 -554 967 -542
rect 932 -571 934 -567
rect 965 -568 967 -564
rect 882 -578 884 -573
rect 891 -587 893 -573
rect 907 -578 909 -573
rect 916 -587 918 -573
rect 78 -596 81 -594
rect 121 -596 139 -594
rect 149 -596 152 -594
rect 34 -621 36 -603
rect 44 -621 46 -603
rect 287 -604 289 -601
rect 297 -604 299 -601
rect 337 -602 339 -599
rect 347 -602 349 -599
rect 78 -606 81 -604
rect 121 -606 139 -604
rect 149 -606 152 -604
rect -27 -637 -25 -625
rect -362 -669 -360 -666
rect -352 -669 -350 -666
rect -300 -667 -298 -663
rect -290 -667 -288 -663
rect -108 -658 -106 -640
rect -98 -658 -96 -640
rect -74 -658 -72 -640
rect -64 -658 -62 -640
rect -9 -641 -7 -623
rect 1 -641 3 -623
rect 253 -624 255 -620
rect 263 -624 265 -620
rect 76 -631 78 -628
rect 86 -631 88 -628
rect -27 -650 -25 -647
rect 34 -645 36 -641
rect 44 -645 46 -641
rect -9 -654 -7 -651
rect 1 -654 3 -651
rect -249 -670 -247 -667
rect -239 -670 -237 -667
rect -396 -680 -394 -676
rect -386 -680 -384 -676
rect -74 -671 -72 -668
rect -64 -671 -62 -668
rect 127 -637 129 -633
rect 137 -637 139 -633
rect 158 -643 160 -639
rect -108 -682 -106 -678
rect -98 -682 -96 -678
rect -880 -710 -878 -698
rect -880 -733 -878 -730
rect -872 -739 -870 -698
rect -856 -710 -854 -698
rect -856 -733 -854 -730
rect -871 -742 -870 -739
rect -848 -742 -846 -698
rect -830 -714 -828 -698
rect -812 -710 -810 -698
rect -803 -710 -801 -706
rect -787 -710 -785 -698
rect -778 -710 -776 -706
rect -830 -728 -828 -724
rect -762 -714 -760 -698
rect -667 -699 -665 -687
rect -658 -699 -656 -696
rect -511 -699 -509 -696
rect -502 -699 -500 -687
rect 76 -689 78 -671
rect 86 -689 88 -671
rect 127 -675 129 -657
rect 137 -675 139 -657
rect 374 -607 376 -603
rect 384 -607 386 -603
rect 464 -607 466 -604
rect 474 -607 476 -604
rect 405 -613 407 -609
rect 253 -662 255 -644
rect 263 -662 265 -644
rect 287 -662 289 -644
rect 297 -662 299 -644
rect 337 -660 339 -642
rect 347 -660 349 -642
rect 374 -645 376 -627
rect 384 -645 386 -627
rect 446 -629 448 -626
rect 405 -645 407 -633
rect 158 -675 160 -663
rect -636 -718 -632 -716
rect -612 -718 -600 -716
rect -590 -718 -586 -716
rect -581 -718 -577 -716
rect -567 -718 -555 -716
rect -535 -718 -531 -716
rect -762 -728 -760 -724
rect -667 -725 -665 -719
rect -812 -735 -810 -730
rect -803 -744 -801 -730
rect -787 -735 -785 -730
rect -778 -744 -776 -730
rect -667 -732 -665 -728
rect -658 -732 -656 -719
rect -454 -705 -452 -693
rect -445 -705 -443 -702
rect -298 -705 -296 -702
rect -289 -705 -287 -693
rect -511 -732 -509 -719
rect -502 -725 -500 -719
rect -423 -724 -419 -722
rect -399 -724 -387 -722
rect -377 -724 -373 -722
rect -368 -724 -364 -722
rect -354 -724 -342 -722
rect -322 -724 -318 -722
rect -502 -732 -500 -728
rect -454 -731 -452 -725
rect -454 -738 -452 -734
rect -445 -738 -443 -725
rect -166 -707 -164 -695
rect -157 -707 -155 -704
rect -10 -707 -8 -704
rect -1 -707 1 -695
rect 812 -608 814 -604
rect 820 -608 822 -604
rect 836 -608 838 -604
rect 844 -608 846 -604
rect 862 -608 864 -604
rect 880 -608 882 -605
rect 905 -608 907 -605
rect 930 -608 932 -604
rect 564 -617 566 -614
rect 574 -617 576 -614
rect 498 -627 500 -623
rect 508 -627 510 -623
rect 529 -633 531 -629
rect 405 -659 407 -655
rect 446 -661 448 -649
rect 374 -669 376 -665
rect 384 -669 386 -665
rect 287 -675 289 -672
rect 297 -675 299 -672
rect 337 -673 339 -670
rect 347 -673 349 -670
rect 464 -665 466 -647
rect 474 -665 476 -647
rect 498 -665 500 -647
rect 508 -665 510 -647
rect 529 -665 531 -653
rect 962 -609 964 -605
rect 592 -639 594 -636
rect 623 -639 625 -635
rect 633 -639 635 -635
rect 446 -674 448 -671
rect 464 -678 466 -675
rect 474 -678 476 -675
rect 158 -689 160 -685
rect 253 -686 255 -682
rect 263 -686 265 -682
rect 564 -675 566 -657
rect 574 -675 576 -657
rect 812 -640 814 -628
rect 592 -671 594 -659
rect 529 -679 531 -675
rect 623 -677 625 -659
rect 633 -677 635 -659
rect 812 -663 814 -660
rect 820 -669 822 -628
rect 836 -640 838 -628
rect 836 -663 838 -660
rect 821 -672 822 -669
rect 844 -672 846 -628
rect 862 -644 864 -628
rect 880 -640 882 -628
rect 889 -640 891 -636
rect 905 -640 907 -628
rect 914 -640 916 -636
rect 862 -658 864 -654
rect 930 -644 932 -628
rect 962 -641 964 -629
rect 930 -658 932 -654
rect 962 -655 964 -651
rect 880 -665 882 -660
rect 889 -674 891 -660
rect 905 -665 907 -660
rect 914 -674 916 -660
rect 592 -684 594 -681
rect 498 -689 500 -685
rect 508 -689 510 -685
rect 564 -688 566 -685
rect 574 -688 576 -685
rect 127 -699 129 -695
rect 137 -699 139 -695
rect 76 -702 78 -699
rect 86 -702 88 -699
rect -298 -738 -296 -725
rect -289 -731 -287 -725
rect -135 -726 -131 -724
rect -111 -726 -99 -724
rect -89 -726 -85 -724
rect -80 -726 -76 -724
rect -66 -726 -54 -724
rect -34 -726 -30 -724
rect -166 -733 -164 -727
rect -289 -738 -287 -734
rect -667 -744 -665 -742
rect -667 -748 -666 -744
rect -658 -745 -656 -742
rect -511 -745 -509 -742
rect -502 -744 -500 -742
rect -501 -748 -500 -744
rect -166 -740 -164 -736
rect -157 -740 -155 -727
rect 195 -711 197 -699
rect 204 -711 206 -708
rect 351 -711 353 -708
rect 360 -711 362 -699
rect 623 -701 625 -697
rect 633 -701 635 -697
rect 808 -700 810 -696
rect 816 -700 818 -696
rect 832 -700 834 -696
rect 840 -700 842 -696
rect 858 -700 860 -696
rect 876 -700 878 -697
rect 901 -700 903 -697
rect 926 -700 928 -696
rect -10 -740 -8 -727
rect -1 -733 1 -727
rect 226 -730 230 -728
rect 250 -730 262 -728
rect 272 -730 276 -728
rect 281 -730 285 -728
rect 295 -730 307 -728
rect 327 -730 331 -728
rect -1 -740 1 -736
rect 195 -737 197 -731
rect -667 -749 -665 -748
rect -502 -749 -500 -748
rect -454 -750 -452 -748
rect -454 -754 -453 -750
rect -445 -751 -443 -748
rect -298 -751 -296 -748
rect -289 -750 -287 -748
rect 195 -744 197 -740
rect 204 -744 206 -731
rect 537 -716 540 -714
rect 580 -716 598 -714
rect 608 -716 611 -714
rect 427 -721 431 -719
rect 451 -721 469 -719
rect 489 -721 493 -719
rect 961 -701 963 -697
rect 537 -726 540 -724
rect 580 -726 598 -724
rect 608 -726 611 -724
rect 427 -731 431 -729
rect 451 -731 469 -729
rect 489 -731 493 -729
rect 351 -744 353 -731
rect 360 -737 362 -731
rect 808 -732 810 -720
rect 360 -744 362 -740
rect -288 -754 -287 -750
rect -454 -755 -452 -754
rect -289 -755 -287 -754
rect -166 -752 -164 -750
rect -166 -756 -165 -752
rect -157 -753 -155 -750
rect -10 -753 -8 -750
rect -1 -752 1 -750
rect 0 -756 1 -752
rect -166 -757 -164 -756
rect -1 -757 1 -756
rect 195 -756 197 -754
rect 195 -760 196 -756
rect 204 -757 206 -754
rect 351 -757 353 -754
rect 360 -756 362 -754
rect 427 -755 431 -753
rect 451 -755 469 -753
rect 489 -755 493 -753
rect 808 -755 810 -752
rect 361 -760 362 -756
rect 195 -761 197 -760
rect 360 -761 362 -760
rect -883 -765 -881 -761
rect -875 -765 -873 -761
rect -859 -765 -857 -761
rect -851 -765 -849 -761
rect -833 -765 -831 -761
rect -815 -765 -813 -762
rect -790 -765 -788 -762
rect -765 -765 -763 -761
rect 816 -761 818 -720
rect 832 -732 834 -720
rect 832 -755 834 -752
rect 427 -765 431 -763
rect 451 -765 469 -763
rect 489 -765 493 -763
rect 817 -764 818 -761
rect 840 -764 842 -720
rect 858 -736 860 -720
rect 876 -732 878 -720
rect 885 -732 887 -728
rect 901 -732 903 -720
rect 910 -732 912 -728
rect 858 -750 860 -746
rect 926 -736 928 -720
rect 961 -733 963 -721
rect 926 -750 928 -746
rect 961 -747 963 -743
rect 876 -757 878 -752
rect 885 -766 887 -752
rect 901 -757 903 -752
rect 910 -766 912 -752
rect -883 -797 -881 -785
rect -883 -820 -881 -817
rect -875 -826 -873 -785
rect -859 -797 -857 -785
rect -859 -820 -857 -817
rect -874 -829 -873 -826
rect -851 -829 -849 -785
rect -833 -801 -831 -785
rect -815 -797 -813 -785
rect -806 -797 -804 -793
rect -790 -797 -788 -785
rect -781 -797 -779 -793
rect -833 -815 -831 -811
rect -765 -801 -763 -785
rect 805 -786 807 -782
rect 813 -786 815 -782
rect 829 -786 831 -782
rect 837 -786 839 -782
rect 855 -786 857 -782
rect 873 -786 875 -783
rect 898 -786 900 -783
rect 923 -786 925 -782
rect 962 -787 964 -783
rect -765 -815 -763 -811
rect -815 -822 -813 -817
rect -806 -831 -804 -817
rect -790 -822 -788 -817
rect -781 -831 -779 -817
rect 805 -818 807 -806
rect 805 -841 807 -838
rect 813 -847 815 -806
rect 829 -818 831 -806
rect 829 -841 831 -838
rect 814 -850 815 -847
rect 837 -850 839 -806
rect 855 -822 857 -806
rect 873 -818 875 -806
rect 882 -818 884 -814
rect 898 -818 900 -806
rect 907 -818 909 -814
rect 855 -836 857 -832
rect 923 -822 925 -806
rect 962 -819 964 -807
rect 923 -836 925 -832
rect 962 -833 964 -829
rect 873 -843 875 -838
rect 882 -852 884 -838
rect 898 -843 900 -838
rect 907 -852 909 -838
rect -882 -862 -880 -858
rect -874 -862 -872 -858
rect -858 -862 -856 -858
rect -850 -862 -848 -858
rect -832 -862 -830 -858
rect -814 -862 -812 -859
rect -789 -862 -787 -859
rect -764 -862 -762 -858
rect -882 -894 -880 -882
rect -882 -917 -880 -914
rect -874 -923 -872 -882
rect -858 -894 -856 -882
rect -858 -917 -856 -914
rect -873 -926 -872 -923
rect -850 -926 -848 -882
rect -832 -898 -830 -882
rect -814 -894 -812 -882
rect -805 -894 -803 -890
rect -789 -894 -787 -882
rect -780 -894 -778 -890
rect -832 -912 -830 -908
rect -764 -898 -762 -882
rect 806 -883 808 -879
rect 814 -883 816 -879
rect 830 -883 832 -879
rect 838 -883 840 -879
rect 856 -883 858 -879
rect 874 -883 876 -880
rect 899 -883 901 -880
rect 924 -883 926 -879
rect 960 -884 962 -880
rect -764 -912 -762 -908
rect -814 -919 -812 -914
rect -805 -928 -803 -914
rect -789 -919 -787 -914
rect -780 -928 -778 -914
rect 806 -915 808 -903
rect 806 -938 808 -935
rect 814 -944 816 -903
rect 830 -915 832 -903
rect 830 -938 832 -935
rect 815 -947 816 -944
rect 838 -947 840 -903
rect 856 -919 858 -903
rect 874 -915 876 -903
rect 883 -915 885 -911
rect 899 -915 901 -903
rect 908 -915 910 -911
rect 856 -933 858 -929
rect 924 -919 926 -903
rect 960 -916 962 -904
rect 924 -933 926 -929
rect 960 -930 962 -926
rect 874 -940 876 -935
rect -884 -952 -882 -948
rect -876 -952 -874 -948
rect -860 -952 -858 -948
rect -852 -952 -850 -948
rect -834 -952 -832 -948
rect -816 -952 -814 -949
rect -791 -952 -789 -949
rect -766 -952 -764 -948
rect 883 -949 885 -935
rect 899 -940 901 -935
rect 908 -949 910 -935
rect -884 -984 -882 -972
rect -884 -1007 -882 -1004
rect -876 -1013 -874 -972
rect -860 -984 -858 -972
rect -860 -1007 -858 -1004
rect -875 -1016 -874 -1013
rect -852 -1016 -850 -972
rect -834 -988 -832 -972
rect -816 -984 -814 -972
rect -807 -984 -805 -980
rect -791 -984 -789 -972
rect -782 -984 -780 -980
rect -834 -1002 -832 -998
rect -766 -988 -764 -972
rect -766 -1002 -764 -998
rect -816 -1009 -814 -1004
rect -807 -1018 -805 -1004
rect -791 -1009 -789 -1004
rect -782 -1018 -780 -1004
rect -885 -1042 -883 -1038
rect -877 -1042 -875 -1038
rect -861 -1042 -859 -1038
rect -853 -1042 -851 -1038
rect -835 -1042 -833 -1038
rect -817 -1042 -815 -1039
rect -792 -1042 -790 -1039
rect -767 -1042 -765 -1038
rect -885 -1074 -883 -1062
rect -885 -1097 -883 -1094
rect -877 -1103 -875 -1062
rect -861 -1074 -859 -1062
rect -861 -1097 -859 -1094
rect -876 -1106 -875 -1103
rect -853 -1106 -851 -1062
rect -835 -1078 -833 -1062
rect -817 -1074 -815 -1062
rect -808 -1074 -806 -1070
rect -792 -1074 -790 -1062
rect -783 -1074 -781 -1070
rect -835 -1092 -833 -1088
rect -767 -1078 -765 -1062
rect -767 -1092 -765 -1088
rect -817 -1099 -815 -1094
rect -808 -1108 -806 -1094
rect -792 -1099 -790 -1094
rect -783 -1108 -781 -1094
rect -886 -1134 -884 -1130
rect -878 -1134 -876 -1130
rect -862 -1134 -860 -1130
rect -854 -1134 -852 -1130
rect -836 -1134 -834 -1130
rect -818 -1134 -816 -1131
rect -793 -1134 -791 -1131
rect -768 -1134 -766 -1130
rect -886 -1166 -884 -1154
rect -886 -1189 -884 -1186
rect -878 -1195 -876 -1154
rect -862 -1166 -860 -1154
rect -862 -1189 -860 -1186
rect -877 -1198 -876 -1195
rect -854 -1198 -852 -1154
rect -836 -1170 -834 -1154
rect -818 -1166 -816 -1154
rect -809 -1166 -807 -1162
rect -793 -1166 -791 -1154
rect -784 -1166 -782 -1162
rect -836 -1184 -834 -1180
rect -768 -1170 -766 -1154
rect -768 -1184 -766 -1180
rect -818 -1191 -816 -1186
rect -809 -1200 -807 -1186
rect -793 -1191 -791 -1186
rect -784 -1200 -782 -1186
rect -884 -1230 -882 -1226
rect -876 -1230 -874 -1226
rect -860 -1230 -858 -1226
rect -852 -1230 -850 -1226
rect -834 -1230 -832 -1226
rect -816 -1230 -814 -1227
rect -791 -1230 -789 -1227
rect -766 -1230 -764 -1226
rect -884 -1262 -882 -1250
rect -884 -1285 -882 -1282
rect -876 -1291 -874 -1250
rect -860 -1262 -858 -1250
rect -860 -1285 -858 -1282
rect -875 -1294 -874 -1291
rect -852 -1294 -850 -1250
rect -834 -1266 -832 -1250
rect -816 -1262 -814 -1250
rect -807 -1262 -805 -1258
rect -791 -1262 -789 -1250
rect -782 -1262 -780 -1258
rect -834 -1280 -832 -1276
rect -766 -1266 -764 -1250
rect -766 -1280 -764 -1276
rect -816 -1287 -814 -1282
rect -807 -1296 -805 -1282
rect -791 -1287 -789 -1282
rect -782 -1296 -780 -1282
<< polycontact >>
rect -878 -531 -874 -527
rect -854 -531 -850 -527
rect -869 -565 -865 -561
rect -846 -565 -842 -561
rect -828 -532 -824 -528
rect -810 -531 -806 -527
rect -785 -531 -781 -527
rect -760 -532 -756 -528
rect -295 -550 -291 -546
rect -801 -565 -797 -561
rect -776 -565 -772 -561
rect -293 -568 -289 -564
rect -299 -578 -295 -574
rect -211 -582 -207 -578
rect -201 -588 -197 -584
rect -880 -618 -876 -614
rect -856 -618 -852 -614
rect -871 -652 -867 -648
rect -848 -652 -844 -648
rect -830 -619 -826 -615
rect -812 -618 -808 -614
rect -787 -618 -783 -614
rect -762 -619 -758 -615
rect -539 -623 -535 -619
rect -803 -652 -799 -648
rect -778 -652 -774 -648
rect -607 -649 -603 -645
rect -597 -643 -593 -639
rect -579 -649 -575 -645
rect -569 -643 -565 -639
rect -515 -649 -511 -645
rect -505 -643 -501 -639
rect -487 -645 -483 -641
rect -466 -645 -462 -641
rect -456 -651 -452 -647
rect -394 -655 -390 -651
rect -384 -649 -380 -645
rect -366 -655 -362 -651
rect -356 -649 -352 -645
rect -319 -642 -315 -638
rect -298 -642 -294 -638
rect -288 -636 -284 -632
rect 810 -552 814 -548
rect -168 -608 -164 -604
rect -158 -602 -154 -598
rect 130 -582 134 -578
rect 834 -552 838 -548
rect -140 -604 -136 -600
rect -247 -650 -243 -646
rect 819 -586 823 -582
rect 842 -586 846 -582
rect 860 -553 864 -549
rect 878 -552 882 -548
rect 903 -552 907 -548
rect 928 -553 932 -549
rect 961 -553 965 -549
rect 887 -586 891 -582
rect 912 -586 916 -582
rect 36 -620 40 -616
rect 128 -600 132 -596
rect 46 -614 50 -610
rect 134 -610 138 -606
rect -25 -636 -21 -632
rect -237 -656 -233 -652
rect -106 -657 -102 -653
rect -96 -651 -92 -647
rect -78 -657 -74 -653
rect -68 -651 -64 -647
rect -7 -634 -3 -630
rect 3 -640 7 -636
rect 123 -668 127 -664
rect -884 -709 -880 -705
rect -860 -709 -856 -705
rect -875 -743 -871 -739
rect -852 -743 -848 -739
rect -834 -710 -830 -706
rect -816 -709 -812 -705
rect -791 -709 -787 -705
rect -766 -710 -762 -706
rect -665 -692 -661 -688
rect -506 -692 -502 -688
rect 72 -688 76 -684
rect 82 -682 86 -678
rect 133 -674 137 -670
rect 370 -638 374 -634
rect 255 -661 259 -657
rect 265 -655 269 -651
rect 283 -661 287 -657
rect 293 -655 297 -651
rect 333 -659 337 -655
rect 343 -653 347 -649
rect 380 -644 384 -640
rect 401 -644 405 -640
rect 154 -674 158 -670
rect -605 -716 -601 -712
rect -566 -716 -562 -712
rect -807 -743 -803 -739
rect -782 -743 -778 -739
rect -452 -698 -448 -694
rect -293 -698 -289 -694
rect -656 -730 -652 -726
rect -515 -730 -511 -726
rect -392 -722 -388 -718
rect -353 -722 -349 -718
rect -164 -700 -160 -696
rect -5 -700 -1 -696
rect 448 -660 452 -656
rect 466 -658 470 -654
rect 494 -657 498 -653
rect 476 -664 480 -660
rect 504 -664 508 -660
rect 525 -664 529 -660
rect 808 -639 812 -635
rect 560 -674 564 -670
rect 570 -668 574 -664
rect 588 -670 592 -666
rect 619 -669 623 -665
rect 629 -676 633 -672
rect 832 -639 836 -635
rect 817 -673 821 -669
rect 840 -673 844 -669
rect 858 -640 862 -636
rect 876 -639 880 -635
rect 901 -639 905 -635
rect 926 -640 930 -636
rect 958 -640 962 -636
rect 885 -673 889 -669
rect 910 -673 914 -669
rect -443 -736 -439 -732
rect -302 -736 -298 -732
rect -104 -724 -100 -720
rect -65 -724 -61 -720
rect -666 -748 -662 -744
rect -505 -748 -501 -744
rect 197 -704 201 -700
rect 356 -704 360 -700
rect -155 -738 -151 -734
rect -14 -738 -10 -734
rect 257 -728 261 -724
rect 296 -728 300 -724
rect -453 -754 -449 -750
rect 593 -714 597 -710
rect 458 -719 462 -715
rect 464 -729 468 -725
rect 587 -724 591 -720
rect 804 -731 808 -727
rect 206 -742 210 -738
rect 347 -742 351 -738
rect -292 -754 -288 -750
rect -165 -756 -161 -752
rect -4 -756 0 -752
rect 458 -753 462 -749
rect 196 -760 200 -756
rect 357 -760 361 -756
rect 464 -763 468 -759
rect 828 -731 832 -727
rect 813 -765 817 -761
rect 836 -765 840 -761
rect 854 -732 858 -728
rect 872 -731 876 -727
rect 897 -731 901 -727
rect 922 -732 926 -728
rect 957 -732 961 -728
rect 881 -765 885 -761
rect 906 -765 910 -761
rect -887 -796 -883 -792
rect -863 -796 -859 -792
rect -878 -830 -874 -826
rect -855 -830 -851 -826
rect -837 -797 -833 -793
rect -819 -796 -815 -792
rect -794 -796 -790 -792
rect -769 -797 -765 -793
rect 801 -817 805 -813
rect -810 -830 -806 -826
rect -785 -830 -781 -826
rect 825 -817 829 -813
rect 810 -851 814 -847
rect 833 -851 837 -847
rect 851 -818 855 -814
rect 869 -817 873 -813
rect 894 -817 898 -813
rect 919 -818 923 -814
rect 958 -818 962 -814
rect 878 -851 882 -847
rect 903 -851 907 -847
rect -886 -893 -882 -889
rect -862 -893 -858 -889
rect -877 -927 -873 -923
rect -854 -927 -850 -923
rect -836 -894 -832 -890
rect -818 -893 -814 -889
rect -793 -893 -789 -889
rect -768 -894 -764 -890
rect 802 -914 806 -910
rect -809 -927 -805 -923
rect -784 -927 -780 -923
rect 826 -914 830 -910
rect 811 -948 815 -944
rect 834 -948 838 -944
rect 852 -915 856 -911
rect 870 -914 874 -910
rect 895 -914 899 -910
rect 920 -915 924 -911
rect 956 -915 960 -911
rect 879 -948 883 -944
rect 904 -948 908 -944
rect -888 -983 -884 -979
rect -864 -983 -860 -979
rect -879 -1017 -875 -1013
rect -856 -1017 -852 -1013
rect -838 -984 -834 -980
rect -820 -983 -816 -979
rect -795 -983 -791 -979
rect -770 -984 -766 -980
rect -811 -1017 -807 -1013
rect -786 -1017 -782 -1013
rect -889 -1073 -885 -1069
rect -865 -1073 -861 -1069
rect -880 -1107 -876 -1103
rect -857 -1107 -853 -1103
rect -839 -1074 -835 -1070
rect -821 -1073 -817 -1069
rect -796 -1073 -792 -1069
rect -771 -1074 -767 -1070
rect -812 -1107 -808 -1103
rect -787 -1107 -783 -1103
rect -890 -1165 -886 -1161
rect -866 -1165 -862 -1161
rect -881 -1199 -877 -1195
rect -858 -1199 -854 -1195
rect -840 -1166 -836 -1162
rect -822 -1165 -818 -1161
rect -797 -1165 -793 -1161
rect -772 -1166 -768 -1162
rect -813 -1199 -809 -1195
rect -788 -1199 -784 -1195
rect -888 -1261 -884 -1257
rect -864 -1261 -860 -1257
rect -879 -1295 -875 -1291
rect -856 -1295 -852 -1291
rect -838 -1262 -834 -1258
rect -820 -1261 -816 -1257
rect -795 -1261 -791 -1257
rect -770 -1262 -766 -1258
rect -811 -1295 -807 -1291
rect -786 -1295 -782 -1291
<< metal1 >>
rect -879 -493 -746 -490
rect -879 -500 -876 -493
rect -855 -500 -852 -493
rect -829 -500 -826 -493
rect -811 -500 -808 -493
rect -786 -500 -783 -493
rect -761 -500 -758 -493
rect 809 -514 942 -511
rect -885 -531 -878 -528
rect -862 -528 -859 -520
rect -870 -531 -854 -528
rect -838 -528 -835 -520
rect -799 -520 -790 -517
rect -774 -520 -765 -517
rect -821 -528 -817 -520
rect -846 -531 -828 -528
rect -870 -532 -867 -531
rect -846 -532 -843 -531
rect -821 -531 -810 -528
rect -793 -528 -790 -520
rect -793 -531 -785 -528
rect -768 -528 -765 -520
rect -753 -528 -749 -520
rect 809 -521 812 -514
rect 833 -521 836 -514
rect 859 -521 862 -514
rect 877 -521 880 -514
rect 902 -521 905 -514
rect 927 -521 930 -514
rect 954 -515 979 -512
rect 960 -522 963 -515
rect -768 -531 -760 -528
rect -821 -536 -817 -531
rect -793 -532 -790 -531
rect -768 -532 -765 -531
rect -753 -531 -687 -528
rect -753 -536 -749 -531
rect -879 -555 -876 -552
rect -855 -555 -852 -552
rect -829 -555 -826 -546
rect -811 -555 -808 -552
rect -786 -555 -783 -552
rect -761 -555 -758 -546
rect -879 -558 -758 -555
rect -885 -565 -869 -562
rect -865 -565 -846 -562
rect -842 -565 -801 -562
rect -797 -565 -776 -562
rect -881 -580 -745 -577
rect -881 -587 -878 -580
rect -857 -587 -854 -580
rect -831 -587 -828 -580
rect -813 -587 -810 -580
rect -788 -587 -785 -580
rect -763 -587 -760 -580
rect -887 -618 -880 -615
rect -864 -615 -861 -607
rect -872 -618 -856 -615
rect -840 -615 -837 -607
rect -801 -607 -792 -604
rect -776 -607 -767 -604
rect -823 -615 -819 -607
rect -848 -618 -830 -615
rect -872 -619 -869 -618
rect -848 -619 -845 -618
rect -823 -618 -812 -615
rect -795 -615 -792 -607
rect -795 -618 -787 -615
rect -770 -615 -767 -607
rect -755 -615 -751 -607
rect -770 -618 -762 -615
rect -823 -623 -819 -618
rect -795 -619 -792 -618
rect -770 -619 -767 -618
rect -755 -618 -703 -615
rect -755 -623 -751 -618
rect -881 -642 -878 -639
rect -857 -642 -854 -639
rect -831 -642 -828 -633
rect -813 -642 -810 -639
rect -788 -642 -785 -639
rect -763 -642 -760 -633
rect -881 -645 -760 -642
rect -887 -652 -871 -649
rect -867 -652 -848 -649
rect -844 -652 -803 -649
rect -799 -652 -778 -649
rect -885 -671 -752 -668
rect -706 -670 -703 -618
rect -690 -662 -687 -531
rect -294 -535 -254 -532
rect -294 -539 -291 -535
rect -296 -542 -284 -539
rect -257 -541 -254 -535
rect -257 -544 -226 -541
rect -213 -544 -138 -541
rect -317 -551 -306 -548
rect -317 -557 -314 -551
rect -294 -557 -291 -550
rect -264 -551 -237 -548
rect -317 -560 -310 -557
rect -317 -575 -314 -560
rect -299 -560 -282 -557
rect -299 -566 -296 -560
rect -300 -569 -296 -566
rect -589 -583 -586 -582
rect -314 -579 -310 -576
rect -581 -583 -485 -582
rect -299 -583 -295 -578
rect -589 -585 -485 -583
rect -589 -602 -586 -585
rect -580 -592 -577 -585
rect -540 -592 -537 -585
rect -516 -592 -513 -585
rect -657 -605 -586 -602
rect -488 -604 -485 -585
rect -376 -589 -373 -588
rect -292 -585 -289 -568
rect -235 -576 -232 -553
rect -242 -579 -232 -576
rect -368 -589 -311 -588
rect -376 -591 -311 -589
rect -235 -589 -232 -579
rect -229 -578 -226 -544
rect -212 -551 -209 -544
rect -194 -551 -190 -544
rect -169 -551 -166 -544
rect -141 -563 -138 -544
rect 753 -552 810 -549
rect 826 -549 829 -541
rect 818 -552 834 -549
rect 850 -549 853 -541
rect 889 -541 898 -538
rect 914 -541 923 -538
rect 867 -549 871 -541
rect 842 -552 860 -549
rect -141 -566 -118 -563
rect -202 -572 -199 -571
rect -202 -575 -190 -572
rect -229 -581 -211 -578
rect -193 -584 -190 -575
rect -141 -573 -138 -566
rect -214 -588 -201 -585
rect -193 -587 -172 -584
rect -121 -585 -118 -566
rect 93 -567 133 -564
rect -23 -576 52 -573
rect 93 -573 96 -567
rect 130 -571 133 -567
rect 65 -576 96 -573
rect 123 -574 135 -571
rect -121 -586 -80 -585
rect -193 -589 -190 -587
rect -614 -612 -610 -605
rect -595 -612 -592 -605
rect -488 -607 -439 -604
rect -531 -619 -528 -612
rect -488 -614 -485 -607
rect -467 -614 -464 -607
rect -449 -614 -445 -607
rect -376 -608 -373 -591
rect -367 -598 -364 -591
rect -314 -595 -311 -591
rect -280 -592 -232 -589
rect -280 -595 -277 -592
rect -317 -598 -277 -595
rect -407 -611 -373 -608
rect -317 -611 -314 -598
rect -305 -605 -301 -598
rect -286 -605 -283 -598
rect -235 -599 -232 -592
rect -175 -598 -172 -587
rect -121 -588 -85 -586
rect -175 -601 -158 -598
rect -150 -600 -147 -591
rect -132 -600 -129 -593
rect -88 -591 -85 -588
rect -80 -591 -51 -590
rect -88 -593 -51 -591
rect -150 -603 -140 -600
rect -172 -607 -168 -604
rect -150 -605 -147 -603
rect -132 -603 -122 -600
rect -132 -605 -129 -603
rect -159 -608 -147 -605
rect -159 -609 -156 -608
rect -401 -618 -397 -611
rect -382 -618 -379 -611
rect -212 -614 -209 -609
rect -88 -610 -85 -593
rect -79 -600 -76 -593
rect -23 -605 -20 -576
rect 5 -583 8 -576
rect 29 -583 33 -576
rect 48 -583 51 -576
rect 38 -604 41 -603
rect 29 -607 41 -604
rect -546 -622 -539 -619
rect -605 -633 -602 -632
rect -614 -636 -602 -633
rect -614 -645 -611 -636
rect -593 -642 -569 -639
rect -561 -641 -558 -632
rect -561 -644 -555 -641
rect -633 -648 -611 -645
rect -614 -650 -611 -648
rect -603 -649 -579 -646
rect -561 -646 -558 -644
rect -570 -649 -558 -646
rect -546 -646 -543 -622
rect -531 -622 -520 -619
rect -221 -617 -173 -614
rect -119 -613 -85 -610
rect -531 -624 -528 -622
rect -540 -639 -537 -634
rect -523 -639 -520 -622
rect -296 -626 -293 -625
rect -540 -642 -527 -639
rect -523 -642 -505 -639
rect -546 -649 -534 -646
rect -588 -650 -583 -649
rect -570 -650 -567 -649
rect -621 -662 -618 -657
rect -690 -665 -618 -662
rect -580 -664 -577 -660
rect -561 -663 -558 -660
rect -885 -678 -882 -671
rect -861 -678 -858 -671
rect -835 -678 -832 -671
rect -817 -678 -814 -671
rect -792 -678 -789 -671
rect -767 -678 -764 -671
rect -706 -674 -701 -670
rect -621 -674 -618 -665
rect -633 -677 -618 -674
rect -595 -675 -592 -670
rect -589 -667 -561 -664
rect -589 -675 -586 -667
rect -747 -683 -646 -680
rect -891 -709 -884 -706
rect -868 -706 -865 -698
rect -876 -709 -860 -706
rect -844 -706 -841 -698
rect -805 -698 -796 -695
rect -780 -698 -771 -695
rect -827 -706 -823 -698
rect -852 -709 -834 -706
rect -876 -710 -873 -709
rect -852 -710 -849 -709
rect -827 -709 -816 -706
rect -799 -706 -796 -698
rect -799 -709 -791 -706
rect -774 -706 -771 -698
rect -759 -706 -755 -698
rect -747 -706 -744 -683
rect -633 -689 -630 -677
rect -595 -678 -586 -675
rect -661 -692 -630 -689
rect -642 -699 -639 -692
rect -774 -709 -766 -706
rect -827 -714 -823 -709
rect -799 -710 -796 -709
rect -774 -710 -771 -709
rect -759 -709 -744 -706
rect -722 -702 -687 -699
rect -759 -714 -755 -709
rect -722 -715 -719 -702
rect -743 -718 -719 -715
rect -885 -733 -882 -730
rect -861 -733 -858 -730
rect -835 -733 -832 -724
rect -817 -733 -814 -730
rect -792 -733 -789 -730
rect -767 -733 -764 -724
rect -885 -736 -764 -733
rect -891 -743 -875 -740
rect -871 -743 -852 -740
rect -848 -743 -807 -740
rect -803 -743 -782 -740
rect -888 -758 -755 -755
rect -888 -765 -885 -758
rect -864 -765 -861 -758
rect -838 -765 -835 -758
rect -820 -765 -817 -758
rect -795 -765 -792 -758
rect -770 -765 -767 -758
rect -894 -796 -887 -793
rect -871 -793 -868 -785
rect -879 -796 -863 -793
rect -847 -793 -844 -785
rect -808 -785 -799 -782
rect -783 -785 -774 -782
rect -830 -793 -826 -785
rect -855 -796 -837 -793
rect -879 -797 -876 -796
rect -855 -797 -852 -796
rect -830 -796 -819 -793
rect -802 -793 -799 -785
rect -802 -796 -794 -793
rect -777 -793 -774 -785
rect -762 -793 -758 -785
rect -743 -793 -740 -718
rect -777 -796 -769 -793
rect -830 -801 -826 -796
rect -802 -797 -799 -796
rect -777 -797 -774 -796
rect -762 -796 -740 -793
rect -733 -733 -695 -730
rect -762 -801 -758 -796
rect -733 -804 -730 -733
rect -698 -746 -695 -733
rect -690 -738 -687 -702
rect -651 -702 -602 -699
rect -585 -702 -582 -686
rect -671 -726 -668 -719
rect -605 -712 -602 -702
rect -587 -706 -580 -702
rect -572 -711 -569 -667
rect -537 -670 -534 -649
rect -530 -662 -527 -642
rect -497 -641 -494 -632
rect -305 -629 -293 -626
rect -479 -641 -476 -634
rect -457 -635 -454 -634
rect -457 -638 -445 -635
rect -497 -644 -487 -641
rect -518 -648 -515 -645
rect -497 -646 -494 -644
rect -479 -644 -466 -641
rect -479 -646 -476 -644
rect -506 -649 -494 -646
rect -506 -650 -503 -649
rect -448 -647 -445 -638
rect -326 -638 -323 -631
rect -305 -638 -302 -629
rect -267 -632 -264 -626
rect -284 -635 -257 -632
rect -392 -639 -389 -638
rect -401 -642 -389 -639
rect -468 -651 -456 -648
rect -448 -650 -439 -647
rect -448 -652 -445 -650
rect -516 -664 -513 -660
rect -497 -664 -494 -660
rect -488 -663 -485 -656
rect -526 -667 -489 -664
rect -442 -668 -439 -650
rect -537 -673 -522 -670
rect -525 -679 -522 -673
rect -442 -671 -426 -668
rect -467 -676 -464 -672
rect -415 -674 -412 -644
rect -401 -651 -398 -642
rect -380 -648 -356 -645
rect -348 -647 -345 -638
rect -329 -641 -323 -638
rect -326 -643 -323 -641
rect -315 -641 -302 -638
rect -305 -643 -302 -641
rect -294 -642 -275 -639
rect -348 -650 -336 -647
rect -260 -648 -257 -635
rect -254 -648 -251 -639
rect -404 -654 -398 -651
rect -401 -656 -398 -654
rect -390 -655 -366 -652
rect -348 -652 -345 -650
rect -357 -655 -345 -652
rect -339 -653 -336 -650
rect -260 -651 -251 -648
rect -243 -649 -230 -646
rect -375 -656 -370 -655
rect -357 -656 -354 -655
rect -521 -683 -481 -680
rect -432 -677 -412 -674
rect -463 -680 -442 -677
rect -432 -685 -429 -677
rect -408 -680 -405 -663
rect -367 -670 -364 -666
rect -348 -668 -345 -666
rect -317 -667 -314 -653
rect -254 -653 -251 -651
rect -254 -656 -242 -653
rect -233 -655 -225 -652
rect -245 -657 -242 -656
rect -348 -670 -318 -668
rect -376 -671 -318 -670
rect -420 -683 -405 -680
rect -382 -681 -379 -676
rect -376 -673 -345 -671
rect -286 -668 -283 -663
rect -313 -671 -277 -668
rect -254 -671 -251 -667
rect -235 -671 -232 -667
rect -221 -671 -218 -617
rect -176 -623 -173 -617
rect -169 -623 -166 -619
rect -150 -623 -147 -619
rect -141 -623 -138 -615
rect -176 -626 -138 -623
rect -113 -620 -109 -613
rect -94 -620 -91 -613
rect 29 -616 32 -607
rect 65 -610 68 -576
rect 50 -613 68 -610
rect 76 -583 103 -580
rect 71 -608 74 -585
rect 130 -589 133 -582
rect 145 -583 156 -580
rect 153 -589 156 -583
rect 121 -592 138 -589
rect 135 -598 138 -592
rect 149 -592 156 -589
rect 71 -611 81 -608
rect 11 -619 32 -616
rect -376 -681 -373 -673
rect -539 -691 -538 -686
rect -533 -689 -532 -686
rect -533 -691 -506 -689
rect -539 -692 -506 -691
rect -420 -686 -417 -683
rect -382 -684 -373 -681
rect -420 -691 -415 -686
rect -539 -693 -532 -692
rect -528 -699 -525 -692
rect -420 -695 -417 -691
rect -448 -698 -417 -695
rect -590 -714 -577 -711
rect -570 -715 -569 -711
rect -565 -702 -516 -699
rect -565 -712 -562 -702
rect -429 -705 -426 -698
rect -438 -708 -389 -705
rect -372 -708 -369 -692
rect -663 -720 -660 -717
rect -612 -723 -600 -720
rect -567 -723 -555 -720
rect -507 -720 -504 -717
rect -680 -728 -668 -726
rect -675 -729 -668 -728
rect -671 -732 -668 -729
rect -663 -732 -660 -725
rect -652 -730 -646 -727
rect -605 -731 -602 -723
rect -635 -734 -602 -731
rect -565 -731 -562 -723
rect -521 -730 -515 -727
rect -565 -734 -532 -731
rect -507 -732 -504 -725
rect -635 -737 -632 -734
rect -535 -737 -532 -734
rect -499 -726 -496 -719
rect -499 -728 -487 -726
rect -499 -729 -492 -728
rect -499 -732 -496 -729
rect -458 -732 -455 -725
rect -392 -718 -389 -708
rect -374 -712 -367 -708
rect -359 -717 -356 -673
rect -281 -674 -218 -671
rect -141 -668 -138 -626
rect -32 -632 -29 -625
rect -14 -632 -11 -623
rect 11 -630 14 -619
rect 29 -621 32 -619
rect 40 -620 54 -617
rect 71 -621 74 -611
rect 128 -617 131 -600
rect 135 -601 139 -598
rect 153 -607 156 -592
rect 273 -595 276 -594
rect 319 -594 366 -592
rect 281 -595 366 -594
rect 273 -597 322 -595
rect 134 -613 138 -610
rect 149 -611 153 -608
rect 71 -624 119 -621
rect 273 -614 276 -597
rect 282 -604 285 -597
rect 332 -602 335 -595
rect 363 -597 366 -595
rect 363 -600 491 -597
rect 369 -607 372 -600
rect 387 -607 391 -600
rect 237 -617 276 -614
rect 400 -613 403 -600
rect -41 -635 -29 -632
rect -104 -641 -101 -640
rect -113 -644 -101 -641
rect -127 -676 -124 -646
rect -113 -651 -110 -644
rect -92 -650 -68 -647
rect -60 -649 -57 -640
rect -41 -643 -38 -635
rect -32 -637 -29 -635
rect -21 -635 -11 -632
rect -3 -633 14 -630
rect 71 -631 74 -624
rect 116 -627 119 -624
rect 237 -627 240 -617
rect 116 -630 240 -627
rect 248 -624 252 -617
rect 267 -624 270 -617
rect 450 -619 453 -600
rect 478 -607 481 -600
rect 439 -622 453 -619
rect 488 -617 491 -600
rect 524 -610 590 -607
rect 524 -617 527 -610
rect 488 -620 527 -617
rect 379 -628 382 -627
rect -14 -637 -11 -635
rect -14 -640 -2 -637
rect 7 -639 11 -636
rect -5 -641 -2 -640
rect 122 -637 125 -630
rect 140 -637 144 -630
rect 48 -646 51 -641
rect 153 -643 156 -630
rect 379 -631 391 -628
rect 450 -629 453 -622
rect 368 -638 370 -634
rect -114 -656 -110 -651
rect -60 -652 -48 -649
rect -113 -658 -110 -656
rect -102 -657 -78 -654
rect -60 -654 -57 -652
rect -69 -657 -57 -654
rect -51 -654 -48 -652
rect -87 -658 -82 -657
rect -69 -658 -66 -657
rect -23 -655 -20 -647
rect -14 -655 -11 -651
rect 5 -655 8 -651
rect 12 -649 60 -646
rect 388 -640 391 -631
rect 493 -627 496 -620
rect 511 -627 515 -620
rect 524 -633 527 -620
rect 559 -617 562 -610
rect 587 -629 590 -610
rect 587 -632 646 -629
rect 409 -640 412 -633
rect 587 -639 590 -632
rect 618 -639 621 -632
rect 636 -639 640 -632
rect 257 -645 260 -644
rect 12 -655 15 -649
rect -23 -658 15 -655
rect -196 -679 -124 -676
rect -312 -685 -309 -683
rect -326 -697 -325 -692
rect -320 -695 -319 -692
rect -196 -694 -193 -679
rect -144 -687 -141 -679
rect -120 -682 -117 -665
rect -79 -672 -76 -668
rect -60 -670 -57 -668
rect -60 -672 -59 -670
rect -132 -685 -117 -682
rect -320 -697 -293 -695
rect -326 -698 -293 -697
rect -262 -697 -193 -694
rect -326 -699 -319 -698
rect -315 -705 -312 -698
rect -377 -720 -364 -717
rect -357 -721 -356 -717
rect -352 -708 -303 -705
rect -352 -718 -349 -708
rect -450 -726 -447 -723
rect -399 -729 -387 -726
rect -354 -729 -342 -726
rect -294 -726 -291 -723
rect -467 -734 -455 -732
rect -690 -741 -678 -738
rect -651 -740 -632 -737
rect -627 -740 -539 -737
rect -535 -739 -519 -737
rect -535 -740 -516 -739
rect -651 -741 -645 -740
rect -698 -749 -686 -746
rect -689 -757 -686 -749
rect -681 -751 -678 -741
rect -648 -745 -645 -741
rect -662 -748 -645 -745
rect -627 -751 -624 -740
rect -681 -754 -624 -751
rect -621 -747 -545 -744
rect -621 -757 -618 -747
rect -689 -760 -618 -757
rect -614 -754 -552 -751
rect -614 -764 -611 -754
rect -725 -767 -611 -764
rect -607 -761 -560 -758
rect -743 -807 -730 -804
rect -888 -820 -885 -817
rect -864 -820 -861 -817
rect -838 -820 -835 -811
rect -820 -820 -817 -817
rect -795 -820 -792 -817
rect -770 -820 -767 -811
rect -888 -823 -767 -820
rect -894 -830 -878 -827
rect -874 -830 -855 -827
rect -851 -830 -810 -827
rect -806 -830 -785 -827
rect -887 -855 -754 -852
rect -887 -862 -884 -855
rect -863 -862 -860 -855
rect -837 -862 -834 -855
rect -819 -862 -816 -855
rect -794 -862 -791 -855
rect -769 -862 -766 -855
rect -893 -893 -886 -890
rect -870 -890 -867 -882
rect -878 -893 -862 -890
rect -846 -890 -843 -882
rect -807 -882 -798 -879
rect -782 -882 -773 -879
rect -829 -890 -825 -882
rect -854 -893 -836 -890
rect -878 -894 -875 -893
rect -854 -894 -851 -893
rect -829 -893 -818 -890
rect -801 -890 -798 -882
rect -801 -893 -793 -890
rect -776 -890 -773 -882
rect -761 -890 -757 -882
rect -743 -890 -740 -807
rect -776 -893 -768 -890
rect -829 -898 -825 -893
rect -801 -894 -798 -893
rect -776 -894 -773 -893
rect -761 -893 -740 -890
rect -761 -898 -757 -893
rect -887 -917 -884 -914
rect -863 -917 -860 -914
rect -837 -917 -834 -908
rect -819 -917 -816 -914
rect -794 -917 -791 -914
rect -769 -917 -766 -908
rect -887 -920 -766 -917
rect -893 -927 -877 -924
rect -873 -927 -854 -924
rect -850 -927 -809 -924
rect -805 -927 -784 -924
rect -889 -945 -756 -942
rect -889 -952 -886 -945
rect -865 -952 -862 -945
rect -839 -952 -836 -945
rect -821 -952 -818 -945
rect -796 -952 -793 -945
rect -771 -952 -768 -945
rect -895 -983 -888 -980
rect -872 -980 -869 -972
rect -880 -983 -864 -980
rect -848 -980 -845 -972
rect -809 -972 -800 -969
rect -784 -972 -775 -969
rect -831 -980 -827 -972
rect -856 -983 -838 -980
rect -880 -984 -877 -983
rect -856 -984 -853 -983
rect -831 -983 -820 -980
rect -803 -980 -800 -972
rect -803 -983 -795 -980
rect -778 -980 -775 -972
rect -763 -980 -759 -972
rect -724 -980 -721 -767
rect -607 -771 -604 -761
rect -778 -983 -770 -980
rect -831 -988 -827 -983
rect -803 -984 -800 -983
rect -778 -984 -775 -983
rect -763 -983 -721 -980
rect -711 -774 -604 -771
rect -601 -767 -567 -764
rect -763 -988 -759 -983
rect -889 -1007 -886 -1004
rect -865 -1007 -862 -1004
rect -839 -1007 -836 -998
rect -821 -1007 -818 -1004
rect -796 -1007 -793 -1004
rect -771 -1007 -768 -998
rect -889 -1010 -768 -1007
rect -895 -1017 -879 -1014
rect -875 -1017 -856 -1014
rect -852 -1017 -811 -1014
rect -807 -1017 -786 -1014
rect -890 -1035 -757 -1032
rect -890 -1042 -887 -1035
rect -866 -1042 -863 -1035
rect -840 -1042 -837 -1035
rect -822 -1042 -819 -1035
rect -797 -1042 -794 -1035
rect -772 -1042 -769 -1035
rect -896 -1073 -889 -1070
rect -873 -1070 -870 -1062
rect -881 -1073 -865 -1070
rect -849 -1070 -846 -1062
rect -810 -1062 -801 -1059
rect -785 -1062 -776 -1059
rect -832 -1070 -828 -1062
rect -857 -1073 -839 -1070
rect -881 -1074 -878 -1073
rect -857 -1074 -854 -1073
rect -832 -1073 -821 -1070
rect -804 -1070 -801 -1062
rect -804 -1073 -796 -1070
rect -779 -1070 -776 -1062
rect -764 -1070 -760 -1062
rect -711 -1070 -708 -774
rect -601 -777 -598 -767
rect -779 -1073 -771 -1070
rect -832 -1078 -828 -1073
rect -804 -1074 -801 -1073
rect -779 -1074 -776 -1073
rect -764 -1073 -708 -1070
rect -701 -780 -598 -777
rect -594 -775 -575 -772
rect -764 -1078 -760 -1073
rect -890 -1097 -887 -1094
rect -866 -1097 -863 -1094
rect -840 -1097 -837 -1088
rect -822 -1097 -819 -1094
rect -797 -1097 -794 -1094
rect -772 -1097 -769 -1088
rect -890 -1100 -769 -1097
rect -896 -1107 -880 -1104
rect -876 -1107 -857 -1104
rect -853 -1107 -812 -1104
rect -808 -1107 -787 -1104
rect -891 -1127 -758 -1124
rect -891 -1134 -888 -1127
rect -867 -1134 -864 -1127
rect -841 -1134 -838 -1127
rect -823 -1134 -820 -1127
rect -798 -1134 -795 -1127
rect -773 -1134 -770 -1127
rect -897 -1165 -890 -1162
rect -874 -1162 -871 -1154
rect -882 -1165 -866 -1162
rect -850 -1162 -847 -1154
rect -811 -1154 -802 -1151
rect -786 -1154 -777 -1151
rect -833 -1162 -829 -1154
rect -858 -1165 -840 -1162
rect -882 -1166 -879 -1165
rect -858 -1166 -855 -1165
rect -833 -1165 -822 -1162
rect -805 -1162 -802 -1154
rect -805 -1165 -797 -1162
rect -780 -1162 -777 -1154
rect -765 -1162 -761 -1154
rect -701 -1162 -698 -780
rect -594 -784 -591 -775
rect -780 -1165 -772 -1162
rect -833 -1170 -829 -1165
rect -805 -1166 -802 -1165
rect -780 -1166 -777 -1165
rect -765 -1165 -698 -1162
rect -687 -787 -591 -784
rect -578 -784 -575 -775
rect -570 -777 -567 -767
rect -563 -771 -560 -761
rect -555 -764 -552 -754
rect -548 -758 -545 -747
rect -542 -752 -539 -740
rect -522 -742 -516 -740
rect -462 -735 -455 -734
rect -458 -738 -455 -735
rect -450 -738 -447 -731
rect -439 -736 -433 -733
rect -392 -737 -389 -729
rect -422 -740 -389 -737
rect -352 -737 -349 -729
rect -308 -736 -302 -733
rect -352 -740 -319 -737
rect -294 -738 -291 -731
rect -522 -745 -519 -742
rect -422 -743 -419 -740
rect -522 -748 -505 -745
rect -435 -745 -419 -743
rect -438 -746 -419 -745
rect -322 -743 -319 -740
rect -286 -732 -283 -725
rect -286 -734 -274 -732
rect -286 -735 -279 -734
rect -286 -738 -283 -735
rect -322 -745 -306 -743
rect -322 -746 -303 -745
rect -438 -748 -432 -746
rect -542 -755 -497 -752
rect -435 -751 -432 -748
rect -449 -754 -432 -751
rect -309 -748 -303 -746
rect -309 -751 -306 -748
rect -309 -754 -292 -751
rect -548 -761 -504 -758
rect -555 -767 -512 -764
rect -563 -774 -519 -771
rect -570 -780 -527 -777
rect -578 -787 -535 -784
rect -765 -1170 -761 -1165
rect -891 -1189 -888 -1186
rect -867 -1189 -864 -1186
rect -841 -1189 -838 -1180
rect -823 -1189 -820 -1186
rect -798 -1189 -795 -1186
rect -773 -1189 -770 -1180
rect -891 -1192 -770 -1189
rect -897 -1199 -881 -1196
rect -877 -1199 -858 -1196
rect -854 -1199 -813 -1196
rect -809 -1199 -788 -1196
rect -889 -1223 -756 -1220
rect -889 -1230 -886 -1223
rect -865 -1230 -862 -1223
rect -839 -1230 -836 -1223
rect -821 -1230 -818 -1223
rect -796 -1230 -793 -1223
rect -771 -1230 -768 -1223
rect -895 -1261 -888 -1258
rect -872 -1258 -869 -1250
rect -880 -1261 -864 -1258
rect -848 -1258 -845 -1250
rect -809 -1250 -800 -1247
rect -784 -1250 -775 -1247
rect -831 -1258 -827 -1250
rect -856 -1261 -838 -1258
rect -880 -1262 -877 -1261
rect -856 -1262 -853 -1261
rect -831 -1261 -820 -1258
rect -803 -1258 -800 -1250
rect -803 -1261 -795 -1258
rect -778 -1258 -775 -1250
rect -763 -1258 -759 -1250
rect -687 -1258 -684 -787
rect -538 -799 -535 -787
rect -530 -792 -527 -780
rect -522 -786 -519 -774
rect -515 -779 -512 -767
rect -507 -771 -504 -761
rect -501 -760 -497 -755
rect -501 -763 -432 -760
rect -262 -760 -259 -697
rect -132 -697 -129 -685
rect -120 -689 -117 -685
rect -94 -683 -91 -678
rect -88 -675 -59 -672
rect -88 -683 -85 -675
rect -94 -686 -85 -683
rect -160 -700 -129 -697
rect -141 -707 -138 -700
rect -150 -710 -101 -707
rect -84 -710 -81 -694
rect -104 -714 -101 -710
rect -170 -734 -167 -727
rect -102 -719 -101 -714
rect -86 -714 -79 -710
rect -71 -719 -68 -675
rect -38 -699 -37 -694
rect -32 -697 -31 -694
rect -32 -699 -5 -697
rect -38 -700 -5 -699
rect -38 -701 -31 -700
rect -27 -707 -24 -700
rect 57 -703 60 -649
rect 248 -648 260 -645
rect 132 -658 135 -657
rect 132 -661 144 -658
rect 96 -667 123 -664
rect 69 -681 82 -678
rect 90 -680 93 -671
rect 96 -680 99 -667
rect 141 -670 144 -661
rect 162 -670 165 -663
rect 120 -674 133 -671
rect 141 -673 154 -670
rect 141 -675 144 -673
rect 162 -673 168 -670
rect 162 -675 165 -673
rect 234 -680 237 -650
rect 248 -655 251 -648
rect 269 -654 293 -651
rect 301 -653 304 -644
rect 312 -652 343 -649
rect 312 -653 315 -652
rect 351 -651 354 -642
rect 363 -644 380 -641
rect 388 -643 401 -640
rect 363 -651 366 -644
rect 388 -645 391 -643
rect 409 -643 421 -640
rect 409 -645 412 -643
rect 247 -660 251 -655
rect 301 -656 315 -653
rect 351 -654 366 -651
rect 248 -662 251 -660
rect 259 -661 283 -658
rect 301 -658 304 -656
rect 292 -661 304 -658
rect 274 -662 279 -661
rect 292 -662 295 -661
rect 308 -663 311 -656
rect 329 -658 333 -655
rect 351 -656 354 -654
rect 342 -659 354 -656
rect 418 -654 421 -643
rect 342 -660 345 -659
rect 90 -683 99 -680
rect 64 -687 72 -684
rect 90 -685 93 -683
rect 81 -688 93 -685
rect 179 -683 237 -680
rect 81 -689 84 -688
rect 71 -703 74 -699
rect 90 -703 93 -699
rect 122 -700 125 -695
rect 153 -699 156 -685
rect 179 -692 182 -683
rect 217 -691 220 -683
rect 241 -686 244 -669
rect 282 -676 285 -672
rect 301 -674 304 -672
rect 369 -670 372 -665
rect 400 -670 403 -655
rect 441 -656 444 -649
rect 459 -656 462 -647
rect 503 -648 506 -647
rect 503 -651 515 -648
rect 434 -659 444 -656
rect 441 -661 444 -659
rect 452 -659 462 -656
rect 470 -657 494 -654
rect 459 -661 462 -659
rect 512 -660 515 -651
rect 533 -660 536 -653
rect 459 -664 471 -661
rect 480 -663 504 -660
rect 512 -663 525 -660
rect 468 -665 471 -664
rect 512 -665 515 -663
rect 533 -665 540 -660
rect 332 -674 335 -670
rect 351 -674 354 -670
rect 363 -673 403 -670
rect 536 -669 540 -665
rect 557 -667 570 -664
rect 578 -666 581 -657
rect 596 -666 599 -659
rect 628 -660 631 -659
rect 628 -663 640 -660
rect 363 -674 366 -673
rect 301 -676 366 -674
rect 273 -677 366 -676
rect 229 -689 244 -686
rect 267 -687 270 -682
rect 273 -679 304 -677
rect 400 -679 403 -673
rect 450 -679 453 -671
rect 459 -679 462 -675
rect 478 -679 481 -675
rect 273 -687 276 -679
rect 164 -695 182 -692
rect 116 -703 152 -700
rect 57 -706 120 -703
rect -104 -720 -101 -719
rect -89 -722 -76 -719
rect -69 -723 -68 -719
rect -64 -710 -15 -707
rect -64 -720 -61 -710
rect -162 -728 -159 -725
rect -111 -731 -99 -728
rect -66 -731 -54 -728
rect -6 -728 -3 -725
rect -179 -736 -167 -734
rect -174 -737 -167 -736
rect -170 -740 -167 -737
rect -162 -740 -159 -733
rect -151 -738 -145 -735
rect -104 -739 -101 -731
rect -134 -742 -101 -739
rect -64 -739 -61 -731
rect -20 -738 -14 -735
rect -64 -742 -31 -739
rect -6 -740 -3 -733
rect -134 -745 -131 -742
rect -147 -747 -131 -745
rect -150 -748 -131 -747
rect -34 -745 -31 -742
rect 2 -734 5 -727
rect 2 -736 14 -734
rect 2 -737 9 -736
rect 2 -740 5 -737
rect -34 -747 -18 -745
rect -34 -748 -15 -747
rect -150 -750 -144 -748
rect -147 -753 -144 -750
rect -161 -756 -144 -753
rect -21 -750 -15 -748
rect -21 -753 -18 -750
rect -21 -756 -4 -753
rect -388 -763 -259 -760
rect -398 -771 -395 -768
rect -507 -774 -395 -771
rect -388 -779 -385 -763
rect -105 -769 -102 -763
rect -515 -782 -385 -779
rect -381 -772 -102 -769
rect -381 -786 -378 -772
rect 164 -775 167 -695
rect 229 -701 232 -689
rect 267 -690 276 -687
rect 201 -704 232 -701
rect 220 -711 223 -704
rect 211 -714 260 -711
rect 277 -714 280 -698
rect 191 -738 194 -731
rect 257 -724 260 -714
rect 275 -718 282 -714
rect 290 -723 293 -679
rect 400 -682 489 -679
rect 337 -692 340 -688
rect 486 -690 489 -682
rect 493 -690 496 -685
rect 524 -689 527 -675
rect 537 -678 540 -669
rect 578 -669 588 -666
rect 552 -672 560 -671
rect 557 -674 560 -672
rect 578 -671 581 -669
rect 596 -669 619 -666
rect 596 -671 599 -669
rect 569 -674 581 -671
rect 569 -675 572 -674
rect 637 -672 640 -663
rect 538 -683 540 -678
rect 618 -676 629 -673
rect 637 -675 650 -672
rect 637 -677 640 -675
rect 559 -689 562 -685
rect 578 -689 581 -685
rect 587 -689 590 -681
rect 524 -690 615 -689
rect 486 -692 615 -690
rect 486 -693 527 -692
rect 323 -703 324 -698
rect 329 -701 330 -698
rect 329 -703 356 -701
rect 323 -704 356 -703
rect 323 -705 330 -704
rect 334 -711 337 -704
rect 272 -726 285 -723
rect 292 -727 293 -723
rect 297 -714 346 -711
rect 297 -724 300 -714
rect 421 -714 424 -708
rect 421 -717 431 -714
rect 199 -732 202 -729
rect 250 -735 262 -732
rect 295 -735 307 -732
rect 355 -732 358 -729
rect 182 -740 194 -738
rect 187 -741 194 -740
rect 191 -744 194 -741
rect 199 -744 202 -737
rect 210 -742 216 -739
rect 257 -743 260 -735
rect 227 -746 260 -743
rect 297 -743 300 -735
rect 341 -742 347 -739
rect 297 -746 330 -743
rect 355 -744 358 -737
rect 227 -749 230 -746
rect 214 -751 230 -749
rect 211 -752 230 -751
rect 327 -749 330 -746
rect 363 -738 366 -731
rect 421 -732 424 -717
rect 458 -715 461 -706
rect 465 -708 468 -700
rect 465 -713 466 -708
rect 451 -727 455 -724
rect 465 -725 468 -713
rect 494 -714 497 -693
rect 489 -717 497 -714
rect 421 -736 431 -732
rect 452 -733 455 -727
rect 452 -736 469 -733
rect 363 -740 375 -738
rect 363 -741 370 -740
rect 363 -744 366 -741
rect 421 -748 424 -736
rect 327 -751 343 -749
rect 327 -752 346 -751
rect 211 -754 217 -752
rect 214 -757 217 -754
rect 200 -760 217 -757
rect 340 -754 346 -752
rect 421 -751 431 -748
rect 340 -757 343 -754
rect 340 -760 357 -757
rect 421 -766 424 -751
rect 458 -749 462 -747
rect 451 -761 455 -758
rect 465 -759 468 -736
rect 494 -748 497 -717
rect 530 -709 533 -707
rect 530 -712 540 -709
rect 530 -737 533 -712
rect 587 -720 590 -695
rect 612 -702 615 -692
rect 647 -695 650 -675
rect 618 -702 621 -697
rect 612 -705 643 -702
rect 593 -710 596 -705
rect 612 -709 615 -705
rect 608 -712 615 -709
rect 753 -712 756 -552
rect 818 -553 821 -552
rect 842 -553 845 -552
rect 867 -552 878 -549
rect 895 -549 898 -541
rect 895 -552 903 -549
rect 920 -549 923 -541
rect 935 -549 939 -541
rect 969 -549 972 -542
rect 920 -552 928 -549
rect 867 -557 871 -552
rect 895 -553 898 -552
rect 920 -553 923 -552
rect 935 -552 961 -549
rect 935 -557 939 -552
rect 969 -552 976 -549
rect 969 -554 972 -552
rect 809 -576 812 -573
rect 833 -576 836 -573
rect 859 -576 862 -567
rect 877 -576 880 -573
rect 902 -576 905 -573
rect 927 -576 930 -567
rect 960 -569 963 -564
rect 954 -572 979 -569
rect 809 -579 930 -576
rect 803 -586 819 -583
rect 823 -586 842 -583
rect 846 -586 887 -583
rect 891 -586 912 -583
rect 807 -601 940 -598
rect 807 -608 810 -601
rect 831 -608 834 -601
rect 857 -608 860 -601
rect 875 -608 878 -601
rect 900 -608 903 -601
rect 925 -608 928 -601
rect 951 -602 976 -599
rect 957 -609 960 -602
rect 594 -722 598 -719
rect 594 -728 597 -722
rect 580 -731 597 -728
rect 612 -728 615 -712
rect 608 -731 615 -728
rect 624 -715 756 -712
rect 761 -639 808 -636
rect 824 -636 827 -628
rect 816 -639 832 -636
rect 848 -636 851 -628
rect 887 -628 896 -625
rect 912 -628 921 -625
rect 865 -636 869 -628
rect 840 -639 858 -636
rect 589 -742 592 -731
rect 624 -736 627 -715
rect 761 -721 764 -639
rect 816 -640 819 -639
rect 840 -640 843 -639
rect 865 -639 876 -636
rect 893 -636 896 -628
rect 893 -639 901 -636
rect 918 -636 921 -628
rect 933 -636 937 -628
rect 966 -636 969 -629
rect 918 -639 926 -636
rect 865 -644 869 -639
rect 893 -640 896 -639
rect 918 -640 921 -639
rect 933 -639 958 -636
rect 933 -644 937 -639
rect 966 -639 973 -636
rect 966 -641 969 -639
rect 807 -663 810 -660
rect 831 -663 834 -660
rect 857 -663 860 -654
rect 875 -663 878 -660
rect 900 -663 903 -660
rect 925 -663 928 -654
rect 957 -656 960 -651
rect 951 -659 976 -656
rect 807 -666 928 -663
rect 801 -673 817 -670
rect 821 -673 840 -670
rect 844 -673 885 -670
rect 889 -673 910 -670
rect 803 -693 936 -690
rect 803 -700 806 -693
rect 827 -700 830 -693
rect 853 -700 856 -693
rect 871 -700 874 -693
rect 896 -700 899 -693
rect 921 -700 924 -693
rect 950 -694 975 -691
rect 956 -701 959 -694
rect 523 -745 592 -742
rect 599 -739 627 -736
rect 632 -724 764 -721
rect 489 -751 497 -748
rect 599 -751 602 -739
rect 632 -743 635 -724
rect -522 -789 -378 -786
rect -374 -778 167 -775
rect -374 -792 -371 -778
rect 244 -783 247 -768
rect 379 -770 382 -766
rect 421 -770 431 -766
rect 452 -767 455 -761
rect 452 -770 469 -767
rect 312 -774 374 -771
rect 379 -773 416 -770
rect 371 -776 374 -774
rect 371 -779 409 -776
rect -530 -795 -371 -792
rect -366 -786 247 -783
rect 287 -783 364 -780
rect 361 -784 364 -783
rect -366 -799 -363 -786
rect 361 -787 401 -784
rect 287 -793 357 -790
rect 354 -795 357 -793
rect 398 -792 401 -787
rect 406 -786 409 -779
rect 413 -780 416 -773
rect 421 -776 424 -770
rect 464 -777 467 -770
rect 494 -773 497 -751
rect 521 -754 602 -751
rect 607 -746 635 -743
rect 639 -731 804 -728
rect 820 -728 823 -720
rect 812 -731 828 -728
rect 844 -728 847 -720
rect 883 -720 892 -717
rect 908 -720 917 -717
rect 861 -728 865 -720
rect 836 -731 854 -728
rect 521 -777 524 -754
rect 607 -759 610 -746
rect 639 -749 642 -731
rect 812 -732 815 -731
rect 836 -732 839 -731
rect 861 -731 872 -728
rect 889 -728 892 -720
rect 889 -731 897 -728
rect 914 -728 917 -720
rect 929 -728 933 -720
rect 965 -728 968 -721
rect 914 -731 922 -728
rect 464 -780 524 -777
rect 530 -762 610 -759
rect 613 -752 642 -749
rect 646 -737 766 -734
rect 861 -736 865 -731
rect 889 -732 892 -731
rect 914 -732 917 -731
rect 929 -731 957 -728
rect 929 -736 933 -731
rect 965 -731 972 -728
rect 965 -733 968 -731
rect 413 -783 459 -780
rect 456 -785 459 -783
rect 530 -785 533 -762
rect 613 -765 616 -752
rect 646 -755 649 -737
rect 406 -789 452 -786
rect 456 -788 533 -785
rect 536 -768 616 -765
rect 619 -758 649 -755
rect 653 -743 758 -740
rect 449 -791 452 -789
rect 536 -791 539 -768
rect 619 -771 622 -758
rect 653 -762 656 -743
rect 398 -795 443 -792
rect 449 -794 539 -791
rect 542 -774 622 -771
rect 626 -765 656 -762
rect 354 -798 394 -795
rect -538 -802 -363 -799
rect 391 -799 394 -798
rect 440 -798 443 -795
rect 542 -798 545 -774
rect 626 -777 629 -765
rect 391 -802 435 -799
rect 440 -801 545 -798
rect 548 -780 629 -777
rect 432 -804 435 -802
rect 548 -804 551 -780
rect 432 -807 551 -804
rect 755 -911 758 -743
rect 763 -814 766 -737
rect 803 -755 806 -752
rect 827 -755 830 -752
rect 853 -755 856 -746
rect 871 -755 874 -752
rect 896 -755 899 -752
rect 921 -755 924 -746
rect 956 -748 959 -743
rect 950 -751 975 -748
rect 803 -758 924 -755
rect 797 -765 813 -762
rect 817 -765 836 -762
rect 840 -765 881 -762
rect 885 -765 906 -762
rect 800 -779 933 -776
rect 800 -786 803 -779
rect 824 -786 827 -779
rect 850 -786 853 -779
rect 868 -786 871 -779
rect 893 -786 896 -779
rect 918 -786 921 -779
rect 951 -780 976 -777
rect 957 -787 960 -780
rect 763 -817 801 -814
rect 817 -814 820 -806
rect 809 -817 825 -814
rect 841 -814 844 -806
rect 880 -806 889 -803
rect 905 -806 914 -803
rect 858 -814 862 -806
rect 833 -817 851 -814
rect 809 -818 812 -817
rect 833 -818 836 -817
rect 858 -817 869 -814
rect 886 -814 889 -806
rect 886 -817 894 -814
rect 911 -814 914 -806
rect 926 -814 930 -806
rect 966 -814 969 -807
rect 911 -817 919 -814
rect 858 -822 862 -817
rect 886 -818 889 -817
rect 911 -818 914 -817
rect 926 -817 958 -814
rect 926 -822 930 -817
rect 966 -817 973 -814
rect 966 -819 969 -817
rect 800 -841 803 -838
rect 824 -841 827 -838
rect 850 -841 853 -832
rect 868 -841 871 -838
rect 893 -841 896 -838
rect 918 -841 921 -832
rect 957 -834 960 -829
rect 951 -837 976 -834
rect 800 -844 921 -841
rect 794 -851 810 -848
rect 814 -851 833 -848
rect 837 -851 878 -848
rect 882 -851 903 -848
rect 801 -876 934 -873
rect 801 -883 804 -876
rect 825 -883 828 -876
rect 851 -883 854 -876
rect 869 -883 872 -876
rect 894 -883 897 -876
rect 919 -883 922 -876
rect 949 -877 974 -874
rect 955 -884 958 -877
rect 755 -914 802 -911
rect 818 -911 821 -903
rect 810 -914 826 -911
rect 842 -911 845 -903
rect 881 -903 890 -900
rect 906 -903 915 -900
rect 859 -911 863 -903
rect 834 -914 852 -911
rect 810 -915 813 -914
rect 834 -915 837 -914
rect 859 -914 870 -911
rect 887 -911 890 -903
rect 887 -914 895 -911
rect 912 -911 915 -903
rect 927 -911 931 -903
rect 964 -911 967 -904
rect 912 -914 920 -911
rect 859 -919 863 -914
rect 887 -915 890 -914
rect 912 -915 915 -914
rect 927 -914 956 -911
rect 927 -919 931 -914
rect 964 -914 971 -911
rect 964 -916 967 -914
rect 801 -938 804 -935
rect 825 -938 828 -935
rect 851 -938 854 -929
rect 869 -938 872 -935
rect 894 -938 897 -935
rect 919 -938 922 -929
rect 955 -931 958 -926
rect 949 -934 974 -931
rect 801 -941 922 -938
rect 795 -948 811 -945
rect 815 -948 834 -945
rect 838 -948 879 -945
rect 883 -948 904 -945
rect -778 -1261 -770 -1258
rect -831 -1266 -827 -1261
rect -803 -1262 -800 -1261
rect -778 -1262 -775 -1261
rect -763 -1261 -684 -1258
rect -763 -1266 -759 -1261
rect -889 -1285 -886 -1282
rect -865 -1285 -862 -1282
rect -839 -1285 -836 -1276
rect -821 -1285 -818 -1282
rect -796 -1285 -793 -1282
rect -771 -1285 -768 -1276
rect -889 -1288 -768 -1285
rect -895 -1295 -879 -1292
rect -875 -1295 -856 -1292
rect -852 -1295 -811 -1292
rect -807 -1295 -786 -1292
<< m2contact >>
rect -218 -544 -213 -539
rect -237 -553 -232 -548
rect -301 -588 -296 -583
rect -292 -590 -287 -585
rect 52 -576 57 -571
rect -629 -638 -623 -633
rect -638 -649 -633 -644
rect -588 -639 -583 -634
rect -555 -645 -550 -640
rect -622 -657 -617 -652
rect -588 -655 -583 -650
rect -701 -675 -696 -670
rect -646 -684 -641 -679
rect -592 -707 -587 -702
rect -580 -707 -575 -702
rect -561 -668 -556 -663
rect -523 -650 -518 -645
rect -415 -644 -410 -639
rect -473 -653 -468 -648
rect -531 -667 -526 -662
rect -489 -668 -484 -663
rect -426 -671 -421 -666
rect -409 -654 -404 -649
rect -375 -645 -370 -640
rect -334 -643 -329 -638
rect -230 -649 -225 -644
rect -409 -663 -404 -658
rect -375 -661 -370 -656
rect -339 -658 -334 -653
rect -526 -684 -521 -679
rect -468 -681 -463 -676
rect -229 -660 -224 -655
rect 71 -585 76 -580
rect -433 -690 -428 -685
rect -664 -725 -659 -720
rect -508 -725 -503 -720
rect -379 -713 -374 -708
rect -367 -713 -362 -708
rect 54 -621 59 -616
rect 126 -622 131 -617
rect -127 -646 -122 -641
rect -141 -673 -136 -668
rect -87 -647 -82 -642
rect 363 -638 368 -633
rect -120 -656 -114 -651
rect -121 -665 -116 -660
rect -87 -663 -82 -658
rect -51 -659 -46 -654
rect -313 -690 -308 -685
rect -145 -692 -140 -687
rect -451 -731 -446 -726
rect -295 -731 -290 -726
rect -432 -764 -427 -759
rect -59 -675 -54 -670
rect -107 -719 -102 -714
rect -91 -715 -86 -710
rect -79 -715 -74 -710
rect -25 -692 -20 -687
rect 234 -650 239 -645
rect 64 -681 69 -676
rect 168 -675 173 -670
rect 274 -651 279 -646
rect 242 -660 247 -655
rect 240 -669 245 -664
rect 274 -667 279 -662
rect 324 -660 329 -655
rect 307 -668 312 -663
rect 63 -692 68 -687
rect 552 -668 557 -663
rect -163 -733 -158 -728
rect -7 -733 -2 -728
rect -106 -763 -101 -758
rect 216 -696 221 -691
rect 270 -719 275 -714
rect 282 -719 287 -714
rect 552 -677 557 -672
rect 533 -683 538 -678
rect 613 -677 618 -672
rect 336 -697 341 -692
rect 420 -708 425 -703
rect 198 -737 203 -732
rect 354 -737 359 -732
rect 466 -713 471 -708
rect 582 -700 587 -695
rect 457 -747 462 -742
rect 378 -766 383 -761
rect 593 -705 598 -700
rect 647 -700 652 -695
rect 518 -745 523 -740
rect 307 -775 312 -770
rect 282 -784 287 -779
rect 282 -794 287 -789
<< pdm12contact >>
rect -632 -715 -627 -710
rect -540 -715 -535 -710
rect -419 -721 -414 -716
rect -327 -721 -322 -716
rect -131 -723 -126 -718
rect -39 -723 -34 -718
rect 230 -727 235 -722
rect 322 -727 327 -722
<< metal2 >>
rect -235 -543 -218 -540
rect -235 -548 -232 -543
rect -383 -579 -360 -576
rect -383 -600 -380 -579
rect -363 -585 -360 -579
rect 57 -575 74 -572
rect 71 -580 74 -575
rect -363 -588 -301 -585
rect -287 -589 -225 -586
rect -472 -603 -380 -600
rect -472 -625 -469 -603
rect -333 -604 -274 -601
rect -637 -628 -469 -625
rect -637 -644 -634 -628
rect -623 -637 -588 -634
rect -629 -654 -626 -638
rect -554 -646 -550 -645
rect -554 -649 -523 -646
rect -657 -657 -626 -654
rect -617 -655 -588 -652
rect -472 -648 -469 -628
rect -423 -650 -420 -617
rect -333 -638 -330 -604
rect -410 -643 -375 -640
rect -228 -644 -225 -589
rect 55 -616 58 -606
rect 64 -621 126 -618
rect 54 -627 57 -621
rect -265 -648 -230 -645
rect -423 -653 -409 -650
rect -629 -669 -626 -657
rect -556 -667 -531 -664
rect -404 -661 -375 -658
rect -265 -654 -262 -648
rect -135 -630 57 -627
rect -225 -648 -180 -645
rect -334 -657 -262 -654
rect -224 -659 -206 -655
rect -484 -667 -468 -664
rect -696 -674 -691 -671
rect -637 -672 -626 -669
rect -637 -680 -634 -672
rect -641 -683 -634 -680
rect -684 -721 -681 -693
rect -684 -724 -664 -721
rect -645 -726 -642 -684
rect -544 -682 -526 -679
rect -471 -680 -468 -667
rect -421 -670 -403 -667
rect -631 -698 -596 -695
rect -631 -710 -628 -698
rect -599 -703 -596 -698
rect -571 -698 -536 -695
rect -599 -706 -592 -703
rect -571 -703 -568 -698
rect -575 -706 -568 -703
rect -539 -710 -536 -698
rect -525 -726 -522 -684
rect -406 -678 -403 -670
rect -406 -681 -309 -678
rect -312 -685 -309 -681
rect -183 -679 -180 -648
rect -135 -652 -132 -630
rect -122 -645 -87 -642
rect -135 -655 -120 -652
rect -116 -663 -87 -660
rect -50 -662 54 -659
rect -136 -673 -59 -670
rect 51 -678 54 -662
rect 64 -676 67 -621
rect 127 -625 318 -622
rect 113 -636 172 -633
rect 169 -670 172 -636
rect 239 -649 274 -646
rect 227 -659 242 -656
rect 227 -676 230 -659
rect 315 -656 318 -625
rect 364 -633 367 -585
rect 315 -659 324 -656
rect 545 -662 548 -637
rect 245 -667 274 -664
rect 545 -663 555 -662
rect 545 -665 552 -663
rect 308 -669 312 -668
rect 308 -672 545 -669
rect 542 -673 545 -672
rect 542 -676 552 -673
rect -183 -682 41 -679
rect 51 -681 64 -678
rect 227 -679 397 -676
rect 609 -676 613 -673
rect -503 -724 -480 -721
rect -483 -805 -480 -724
rect -471 -727 -468 -699
rect -471 -730 -451 -727
rect -432 -732 -429 -690
rect -308 -689 -241 -686
rect -418 -704 -383 -701
rect -418 -716 -415 -704
rect -386 -709 -383 -704
rect -358 -704 -323 -701
rect -386 -712 -379 -709
rect -358 -709 -355 -704
rect -362 -712 -355 -709
rect -326 -716 -323 -704
rect -312 -732 -309 -690
rect -290 -730 -267 -727
rect -431 -759 -428 -737
rect -270 -779 -267 -730
rect -183 -729 -180 -701
rect -183 -732 -163 -729
rect -144 -734 -141 -692
rect 38 -688 41 -682
rect 38 -691 63 -688
rect -130 -706 -95 -703
rect -130 -718 -127 -706
rect -98 -711 -95 -706
rect -70 -706 -35 -703
rect -98 -714 -91 -711
rect -70 -711 -67 -706
rect -74 -714 -67 -711
rect -38 -718 -35 -706
rect -106 -758 -103 -719
rect -24 -734 -21 -692
rect -2 -732 21 -729
rect 18 -771 21 -732
rect 178 -733 181 -705
rect 178 -736 198 -733
rect 217 -738 220 -696
rect 394 -694 397 -679
rect 394 -697 404 -694
rect 231 -710 266 -707
rect 231 -722 234 -710
rect 263 -715 266 -710
rect 291 -710 326 -707
rect 263 -718 270 -715
rect 291 -715 294 -710
rect 287 -718 294 -715
rect 323 -722 326 -710
rect 337 -738 340 -697
rect 534 -694 537 -683
rect 534 -695 587 -694
rect 534 -697 582 -695
rect 593 -699 647 -696
rect 593 -700 598 -699
rect 425 -707 429 -704
rect 517 -706 528 -703
rect 471 -713 507 -710
rect 504 -728 507 -713
rect 359 -736 382 -733
rect 379 -761 382 -736
rect 458 -742 518 -741
rect 462 -744 518 -742
rect 18 -772 176 -771
rect 18 -774 307 -772
rect 173 -775 307 -774
rect -270 -782 282 -779
rect -360 -792 282 -789
rect -360 -805 -357 -792
rect -483 -808 -357 -805
<< m3contact >>
rect -424 -617 -419 -612
rect -554 -654 -549 -649
rect -274 -605 -269 -600
rect -206 -660 -201 -655
rect -685 -693 -680 -688
rect 108 -637 113 -632
rect -472 -699 -467 -694
rect -241 -690 -236 -685
rect -184 -701 -179 -696
rect 177 -705 182 -700
rect 404 -698 409 -693
<< m123contact >>
rect -586 -583 -581 -578
rect -373 -589 -368 -584
rect -319 -580 -314 -575
rect -219 -589 -214 -584
rect -268 -626 -263 -621
rect -275 -643 -270 -638
rect -85 -591 -80 -586
rect 276 -595 281 -590
rect -177 -609 -172 -604
rect 153 -612 158 -607
rect -586 -686 -581 -681
rect -538 -691 -533 -686
rect -318 -672 -313 -667
rect 11 -641 16 -636
rect -42 -648 -37 -643
rect 135 -618 140 -613
rect 115 -675 120 -670
rect 434 -622 439 -617
rect 417 -659 422 -654
rect -680 -733 -675 -728
rect -646 -731 -641 -726
rect -526 -731 -521 -726
rect -492 -733 -487 -728
rect -415 -691 -410 -686
rect -373 -692 -368 -687
rect -325 -697 -320 -692
rect -467 -739 -462 -734
rect -433 -737 -428 -732
rect -313 -737 -308 -732
rect -279 -739 -274 -734
rect -399 -768 -394 -763
rect -85 -694 -80 -689
rect 336 -688 341 -683
rect -37 -699 -32 -694
rect -179 -741 -174 -736
rect -145 -739 -140 -734
rect 152 -704 157 -699
rect -25 -739 -20 -734
rect 9 -741 14 -736
rect 232 -697 237 -692
rect 276 -698 281 -693
rect 324 -703 329 -698
rect 457 -706 462 -701
rect 528 -707 533 -702
rect 182 -745 187 -740
rect 216 -743 221 -738
rect 336 -743 341 -738
rect 370 -745 375 -740
rect 243 -768 248 -763
<< metal3 >>
rect -328 -571 -219 -568
rect -388 -575 -355 -572
rect -585 -681 -582 -583
rect -388 -595 -385 -575
rect -358 -580 -355 -575
rect -328 -580 -325 -571
rect -358 -583 -325 -580
rect -423 -598 -385 -595
rect -423 -611 -420 -598
rect -425 -612 -418 -611
rect -425 -617 -424 -612
rect -419 -617 -418 -612
rect -425 -618 -418 -617
rect -555 -649 -548 -648
rect -555 -654 -554 -649
rect -549 -654 -548 -649
rect -555 -655 -548 -654
rect -554 -671 -550 -655
rect -430 -671 -426 -637
rect -554 -675 -426 -671
rect -686 -688 -679 -687
rect -686 -693 -685 -688
rect -680 -690 -679 -688
rect -539 -690 -538 -686
rect -680 -691 -538 -690
rect -533 -691 -532 -686
rect -410 -690 -406 -687
rect -372 -687 -369 -589
rect -318 -667 -315 -580
rect -222 -588 -219 -571
rect -95 -581 -72 -578
rect -218 -593 -215 -589
rect -95 -593 -92 -581
rect -75 -585 -72 -581
rect -75 -588 126 -585
rect -218 -596 -92 -593
rect -275 -600 -268 -599
rect -275 -605 -274 -600
rect -269 -601 -268 -600
rect -269 -604 -176 -601
rect -269 -605 -268 -604
rect -275 -606 -268 -605
rect -179 -607 -177 -604
rect -268 -621 -263 -618
rect -680 -693 -532 -691
rect -686 -694 -679 -693
rect -473 -694 -466 -693
rect -473 -699 -472 -694
rect -467 -696 -466 -694
rect -326 -696 -325 -692
rect -467 -697 -325 -696
rect -320 -697 -319 -692
rect -467 -699 -319 -697
rect -473 -700 -466 -699
rect -274 -713 -271 -643
rect -206 -654 -202 -637
rect -207 -655 -200 -654
rect -207 -660 -206 -655
rect -201 -660 -200 -655
rect -207 -661 -200 -660
rect -242 -685 -235 -684
rect -242 -690 -241 -685
rect -236 -688 -168 -685
rect -236 -690 -235 -688
rect -84 -689 -81 -591
rect 123 -613 126 -588
rect 123 -616 135 -613
rect 107 -632 114 -631
rect 107 -633 108 -632
rect 15 -636 108 -633
rect 16 -639 18 -636
rect 107 -637 108 -636
rect 113 -637 114 -632
rect 107 -638 114 -637
rect -41 -666 -38 -648
rect -41 -669 -25 -666
rect 105 -674 115 -671
rect -242 -691 -235 -690
rect -185 -696 -178 -695
rect -185 -701 -184 -696
rect -179 -698 -178 -696
rect -38 -698 -37 -694
rect -179 -699 -37 -698
rect -32 -699 -31 -694
rect 105 -695 108 -674
rect 44 -698 108 -695
rect 154 -699 157 -612
rect 237 -693 248 -692
rect 277 -693 280 -595
rect 418 -682 421 -659
rect 435 -675 438 -622
rect 435 -678 449 -675
rect 317 -688 336 -685
rect 418 -685 440 -682
rect 403 -693 410 -692
rect 237 -695 243 -693
rect 403 -698 404 -693
rect 409 -696 417 -693
rect 409 -698 410 -696
rect -179 -701 -31 -699
rect -185 -702 -178 -701
rect 176 -700 183 -699
rect 176 -705 177 -700
rect 182 -702 183 -700
rect 323 -702 324 -698
rect 182 -703 324 -702
rect 329 -703 330 -698
rect 403 -699 410 -698
rect 437 -697 440 -685
rect 446 -684 449 -678
rect 446 -687 485 -684
rect 482 -695 485 -687
rect 437 -700 461 -697
rect 482 -698 532 -695
rect 182 -705 330 -703
rect 457 -701 461 -700
rect 176 -706 183 -705
rect 529 -702 532 -698
rect -409 -716 -271 -713
rect -678 -728 -646 -727
rect -675 -730 -646 -728
rect -521 -728 -489 -727
rect -521 -730 -492 -728
rect -491 -746 -488 -733
rect -465 -734 -433 -733
rect -462 -736 -433 -734
rect -409 -746 -406 -716
rect -308 -734 -276 -733
rect -308 -736 -279 -734
rect -177 -736 -145 -735
rect -174 -738 -145 -736
rect -20 -736 12 -735
rect -20 -738 9 -736
rect 184 -740 216 -739
rect 187 -742 216 -740
rect 341 -740 373 -739
rect 341 -742 370 -740
rect -491 -749 -406 -746
rect -398 -763 -395 -759
rect 244 -763 247 -759
<< m234contact >>
rect -691 -675 -686 -670
rect -549 -684 -544 -679
rect -485 -685 -480 -680
rect 363 -585 368 -580
rect 54 -606 59 -601
rect 544 -637 549 -632
rect 604 -677 609 -672
rect 429 -709 434 -704
rect 512 -708 517 -703
rect 503 -733 508 -728
<< m4contact >>
rect -430 -637 -425 -632
rect -268 -618 -263 -613
rect -206 -637 -201 -632
rect -168 -688 -163 -683
rect -25 -669 -20 -664
rect 39 -699 44 -694
rect 312 -689 317 -684
rect 417 -696 422 -691
<< metal4 >>
rect -267 -557 -112 -554
rect -267 -613 -264 -557
rect -115 -564 -112 -557
rect 83 -557 150 -554
rect 83 -564 86 -557
rect -115 -567 86 -564
rect 147 -569 150 -557
rect 147 -572 166 -569
rect 163 -598 166 -572
rect 262 -584 363 -581
rect 262 -598 265 -584
rect 163 -601 265 -598
rect 424 -597 548 -594
rect 59 -605 109 -602
rect -425 -637 -206 -633
rect 106 -649 109 -605
rect 424 -649 427 -597
rect 545 -632 548 -597
rect 106 -652 427 -649
rect -20 -668 214 -665
rect -686 -674 -621 -671
rect -624 -680 -621 -674
rect -624 -683 -549 -680
rect -484 -753 -481 -685
rect -163 -687 32 -684
rect 29 -696 32 -687
rect 211 -686 214 -668
rect 211 -689 312 -686
rect 29 -699 39 -696
rect 605 -692 608 -677
rect 422 -695 608 -692
rect 434 -707 512 -704
rect 107 -715 393 -712
rect 107 -737 110 -715
rect -385 -740 110 -737
rect -385 -742 -382 -740
rect -413 -745 -382 -742
rect -413 -753 -410 -745
rect -484 -756 -410 -753
rect 390 -757 393 -715
rect 504 -757 507 -733
rect 390 -760 507 -757
<< m345contact >>
rect -406 -691 -401 -686
rect 243 -698 248 -693
rect -399 -759 -394 -754
rect 243 -759 248 -754
<< metal5 >>
rect -401 -691 -395 -687
rect -398 -754 -395 -691
rect 244 -754 247 -698
<< labels >>
rlabel metal1 -584 -704 -584 -704 3 vdd
rlabel metal1 -584 -712 -584 -712 3 gnd
rlabel metal1 -598 -604 -598 -604 5 vdd
rlabel metal1 -569 -665 -569 -665 1 gnd
rlabel metal1 -579 -584 -579 -583 5 vdd
rlabel metal1 -445 -650 -439 -647 7 c1
rlabel metal1 -452 -679 -452 -679 1 gnd
rlabel metal1 -461 -606 -461 -606 5 vdd
rlabel m2contact -522 -647 -518 -646 1 p0_inv
rlabel metal1 -478 -643 -476 -640 1 temp100
rlabel metal1 -515 -584 -515 -583 5 vdd
rlabel metal1 -505 -665 -505 -665 1 gnd
rlabel metal1 -530 -621 -528 -618 1 c0_inv
rlabel metal1 -545 -622 -543 -620 3 c0
rlabel metal1 -539 -641 -539 -641 1 gnd
rlabel metal1 -540 -583 -540 -583 5 vdd
rlabel metal2 -482 -750 -481 -748 1 s0
rlabel metal2 -683 -723 -679 -721 3 mid_s0
rlabel metal1 -591 -642 -580 -639 1 a0
rlabel metal1 -591 -649 -580 -646 1 b0
rlabel metal1 -620 -648 -614 -645 1 g0_inv
rlabel metal1 -558 -644 -553 -641 1 p0_inv
rlabel m2contact -472 -651 -468 -649 1 g0_inv
rlabel metal1 -371 -710 -371 -710 3 vdd
rlabel metal1 -371 -718 -371 -718 3 gnd
rlabel metal1 -385 -610 -385 -610 5 vdd
rlabel metal1 -356 -671 -356 -671 1 gnd
rlabel metal1 -366 -590 -366 -589 5 vdd
rlabel metal2 -470 -728 -470 -728 1 mid_s1
rlabel metal2 -269 -756 -268 -754 8 s1
rlabel metal1 -407 -654 -401 -651 1 g1_inv
rlabel metal1 -345 -650 -340 -647 1 p1_inv
rlabel metal1 -378 -648 -367 -645 1 a1
rlabel metal1 -378 -655 -367 -652 1 b1
rlabel metal1 -311 -686 -309 -683 1 c1
rlabel metal1 -233 -591 -233 -590 5 vdd
rlabel metal1 -243 -672 -243 -672 1 gnd
rlabel metal1 -232 -649 -228 -647 7 p1_inv
rlabel metal1 -231 -655 -226 -653 7 p0_inv
rlabel metal1 -259 -651 -255 -649 3 temp101
rlabel metal1 -289 -597 -289 -597 5 vdd
rlabel metal1 -298 -670 -298 -670 1 gnd
rlabel metal1 -282 -641 -278 -640 1 c0
rlabel metal1 -326 -640 -324 -638 1 temp102
rlabel metal1 -315 -568 -315 -568 3 gnd
rlabel metal1 -234 -578 -233 -578 7 vdd
rlabel space -298 -584 -295 -581 1 g0_inv
rlabel metal1 -293 -542 -290 -539 1 temp103
rlabel metal1 -206 -543 -206 -543 5 vdd
rlabel metal1 -197 -616 -197 -616 1 gnd
rlabel metal1 -190 -587 -184 -584 7 temp104
rlabel metal1 -168 -543 -168 -542 5 vdd
rlabel metal1 -158 -624 -158 -624 1 gnd
rlabel metal1 -131 -602 -129 -600 1 c2
rlabel m123contact -218 -587 -218 -587 1 g1_inv
rlabel metal1 -83 -712 -83 -712 3 vdd
rlabel metal1 -83 -720 -83 -720 3 gnd
rlabel metal1 -97 -612 -97 -612 5 vdd
rlabel metal1 -68 -673 -68 -673 1 gnd
rlabel metal1 -78 -592 -78 -591 5 vdd
rlabel metal2 -181 -731 -180 -729 1 mid_s2
rlabel metal2 19 -758 21 -756 8 s2
rlabel metal1 -90 -650 -79 -647 1 a2
rlabel metal1 -90 -657 -79 -654 1 b2
rlabel metal1 -57 -652 -52 -649 1 p2_inv
rlabel metal1 52 -620 54 -618 1 g2_inv
rlabel metal1 65 -687 70 -685 1 p1_inv
rlabel metal1 129 -574 132 -571 1 temp107
rlabel metal1 67 -681 71 -679 1 p2_inv
rlabel metal1 94 -683 98 -681 1 temp105
rlabel metal1 117 -673 121 -672 1 c1
rlabel metal1 163 -672 165 -670 1 temp106
rlabel metal1 23 -619 29 -616 1 temp108
rlabel metal1 -32 -634 -30 -632 1 c3
rlabel metal1 -3 -656 -3 -656 1 gnd
rlabel metal1 7 -575 7 -574 5 vdd
rlabel metal1 36 -648 36 -648 1 gnd
rlabel metal1 45 -575 45 -575 5 vdd
rlabel metal1 72 -610 73 -610 3 vdd
rlabel metal1 154 -600 154 -600 7 gnd
rlabel metal1 137 -702 137 -702 1 gnd
rlabel metal1 128 -629 128 -629 5 vdd
rlabel metal1 82 -704 82 -704 1 gnd
rlabel metal1 72 -623 72 -622 5 vdd
rlabel m2contact -22 -690 -22 -690 1 c2
rlabel m2contact -120 -655 -114 -652 1 g2_inv
rlabel metal1 135 -616 138 -613 1 g1_inv
rlabel metal1 283 -596 283 -595 5 vdd
rlabel metal1 293 -677 293 -677 1 gnd
rlabel metal1 264 -616 264 -616 5 vdd
rlabel metal1 278 -724 278 -724 3 gnd
rlabel metal1 278 -716 278 -716 3 vdd
rlabel metal2 179 -735 179 -735 1 mid_s3
rlabel metal2 380 -762 382 -760 8 s3
rlabel metal1 338 -697 339 -690 1 c3
rlabel metal1 271 -661 282 -658 1 b3
rlabel metal1 271 -654 282 -651 1 a3
rlabel metal1 242 -660 248 -657 1 g3_inv
rlabel metal1 304 -656 309 -653 1 p3_inv
rlabel metal1 333 -594 333 -593 5 vdd
rlabel metal1 343 -675 343 -675 1 gnd
rlabel metal1 328 -652 332 -650 3 p3_inv
rlabel m2contact 327 -657 329 -656 3 p2_inv
rlabel metal1 357 -654 358 -652 7 temp109
rlabel metal1 375 -599 375 -599 5 vdd
rlabel metal1 384 -672 384 -672 1 gnd
rlabel m2contact 365 -637 368 -634 1 temp101
rlabel metal1 410 -642 412 -640 1 p4
rlabel metal1 499 -619 499 -619 5 vdd
rlabel metal1 508 -692 508 -692 1 gnd
rlabel metal1 535 -662 535 -660 1 temp110
rlabel metal1 470 -680 470 -680 1 gnd
rlabel metal1 480 -599 480 -598 5 vdd
rlabel metal1 487 -662 487 -662 1 temp109
rlabel metal1 481 -657 493 -654 1 temp104
rlabel metal1 441 -658 441 -658 1 temp110
rlabel metal1 560 -609 560 -608 5 vdd
rlabel metal1 570 -690 570 -690 1 gnd
rlabel metal1 597 -668 599 -666 1 temp111
rlabel m2contact 554 -667 557 -665 1 g2_inv
rlabel m2contact 556 -674 556 -674 1 p3_inv
rlabel metal1 624 -631 624 -631 5 vdd
rlabel metal1 633 -704 633 -704 1 gnd
rlabel metal1 640 -675 646 -672 7 temp112
rlabel metal1 531 -710 532 -710 3 vdd
rlabel metal1 613 -720 613 -720 7 gnd
rlabel metal1 590 -736 592 -733 1 g4_inv
rlabel m2contact 615 -676 617 -673 1 g3_inv
rlabel metal1 423 -720 423 -720 3 vdd
rlabel metal1 496 -729 496 -729 7 gnd
rlabel metal1 458 -713 461 -711 5 p4
rlabel metal1 423 -754 423 -754 3 vdd
rlabel metal1 496 -763 496 -763 7 gnd
rlabel metal1 466 -748 467 -746 7 temp113
rlabel m2contact 458 -747 461 -744 7 g4_inv
rlabel metal1 464 -776 467 -770 1 c4
rlabel m2contact 467 -713 470 -710 5 c0
rlabel metal1 -685 -663 -685 -663 3 b0
rlabel metal1 -687 -681 -687 -681 3 a0
rlabel metal1 -719 -701 -719 -701 3 a1
rlabel metal1 -721 -733 -718 -730 3 b1
rlabel metal1 -725 -767 -722 -764 3 a2
rlabel m2contact -524 -681 -523 -681 1 c0
rlabel metal1 -705 -672 -705 -672 1 c0
rlabel metal1 709 -713 709 -713 1 c4
rlabel metal1 707 -723 711 -721 1 s3
rlabel metal1 709 -729 709 -729 1 s2
rlabel metal1 708 -735 708 -735 1 s1
rlabel metal1 708 -741 708 -741 1 s0
rlabel metal1 -878 -492 -878 -492 5 vdd
rlabel metal1 -883 -564 -883 -564 1 clk
rlabel metal1 -860 -557 -860 -557 1 gnd
rlabel metal1 -862 -644 -862 -644 1 gnd
rlabel metal1 -885 -651 -885 -651 1 clk
rlabel metal1 -880 -579 -880 -579 5 vdd
rlabel metal1 -884 -670 -884 -670 5 vdd
rlabel metal1 -889 -742 -889 -742 1 clk
rlabel metal1 -866 -735 -866 -735 1 gnd
rlabel metal1 -887 -757 -887 -757 5 vdd
rlabel metal1 -892 -829 -892 -829 1 clk
rlabel metal1 -869 -822 -869 -822 1 gnd
rlabel metal1 -886 -854 -886 -854 5 vdd
rlabel metal1 -891 -926 -891 -926 1 clk
rlabel metal1 -868 -919 -868 -919 1 gnd
rlabel metal1 -888 -944 -888 -944 5 vdd
rlabel metal1 -893 -1016 -893 -1016 1 clk
rlabel metal1 -870 -1009 -870 -1009 1 gnd
rlabel metal1 -889 -1034 -889 -1034 5 vdd
rlabel metal1 -894 -1106 -894 -1106 1 clk
rlabel metal1 -871 -1099 -871 -1099 1 gnd
rlabel metal1 -890 -1126 -890 -1126 5 vdd
rlabel metal1 -895 -1198 -895 -1198 1 clk
rlabel metal1 -872 -1191 -872 -1191 1 gnd
rlabel metal1 810 -513 810 -513 5 vdd
rlabel metal1 805 -585 805 -585 1 clk
rlabel metal1 828 -578 828 -578 1 gnd
rlabel metal1 826 -665 826 -665 1 gnd
rlabel metal1 803 -672 803 -672 1 clk
rlabel metal1 808 -600 808 -600 5 vdd
rlabel metal1 801 -778 801 -778 5 vdd
rlabel metal1 796 -850 796 -850 1 clk
rlabel metal1 819 -843 819 -843 1 gnd
rlabel metal1 802 -875 802 -875 5 vdd
rlabel metal1 797 -947 797 -947 1 clk
rlabel metal1 820 -940 820 -940 1 gnd
rlabel metal1 -693 -773 -693 -773 1 b2
rlabel metal1 -650 -778 -650 -778 1 a3
rlabel metal1 -620 -785 -620 -785 1 b3
rlabel metal1 -888 -1222 -888 -1222 5 vdd
rlabel metal1 -893 -1294 -893 -1294 1 clk
rlabel metal1 -870 -1287 -870 -1287 1 gnd
rlabel metal1 -885 -530 -883 -528 1 b0_in
rlabel metal1 -886 -617 -886 -617 1 c0_in
rlabel metal1 -889 -707 -889 -707 1 a0_in
rlabel metal1 -893 -892 -891 -890 3 b1_in
rlabel metal1 -895 -983 -893 -980 3 a2_in
rlabel metal1 -896 -1073 -893 -1070 3 b2_in
rlabel metal1 -897 -1164 -895 -1162 3 a3_in
rlabel metal1 938 -552 940 -550 1 c4_out
rlabel metal1 937 -639 939 -637 1 s3_out
rlabel metal1 929 -817 932 -814 1 s1_out
rlabel metal1 930 -914 934 -912 1 s0_out
rlabel metal1 804 -692 804 -692 5 vdd
rlabel metal1 799 -764 799 -764 1 clk
rlabel metal1 822 -757 822 -757 1 gnd
rlabel metal1 932 -731 935 -729 1 s2_out
rlabel metal1 960 -513 960 -513 5 vdd
rlabel metal1 961 -571 961 -571 1 gnd
rlabel metal1 957 -600 957 -600 5 vdd
rlabel metal1 958 -658 958 -658 1 gnd
rlabel metal1 969 -551 972 -549 1 c4_inv
rlabel metal1 957 -778 957 -778 5 vdd
rlabel metal1 958 -836 958 -836 1 gnd
rlabel metal1 967 -638 969 -636 1 s3_inv
rlabel metal1 956 -692 956 -692 5 vdd
rlabel metal1 957 -750 957 -750 1 gnd
rlabel metal1 965 -730 968 -728 1 s2_inv
rlabel metal1 966 -816 969 -814 1 s1_inv
rlabel metal1 955 -875 955 -875 5 vdd
rlabel metal1 956 -933 956 -933 1 gnd
rlabel metal1 964 -913 967 -911 1 s0_inv
rlabel metal1 -894 -795 -892 -793 3 a1_in
rlabel metal1 -895 -1261 -892 -1258 3 b3_in
<< end >>
