magic
tech scmos
timestamp 1731407297
<< nwell >>
rect -3 -138 31 -118
rect -37 -170 31 -138
rect 37 -140 95 -118
rect 37 -150 144 -140
rect 61 -170 144 -150
rect 89 -172 144 -170
rect -95 -257 -62 -225
rect -55 -262 -23 -236
rect 22 -262 54 -236
rect 61 -257 94 -225
<< ntransistor >>
rect 48 -166 50 -156
rect -26 -202 -24 -182
rect -16 -202 -14 -182
rect 8 -192 10 -182
rect 18 -192 20 -182
rect 72 -192 74 -182
rect 82 -192 84 -182
rect 100 -188 102 -178
rect 121 -204 123 -184
rect 131 -204 133 -184
rect -17 -250 -7 -248
rect 6 -250 16 -248
rect -84 -274 -82 -264
rect -75 -274 -73 -264
rect 72 -274 74 -264
rect 81 -274 83 -264
<< ptransistor >>
rect -26 -164 -24 -144
rect -16 -164 -14 -144
rect 8 -164 10 -124
rect 18 -164 20 -124
rect 48 -144 50 -124
rect 72 -164 74 -124
rect 82 -164 84 -124
rect 100 -166 102 -146
rect 121 -166 123 -146
rect 131 -166 133 -146
rect -84 -251 -82 -231
rect -75 -251 -73 -231
rect -49 -250 -29 -248
rect 28 -250 48 -248
rect 72 -251 74 -231
rect 81 -251 83 -231
<< ndiffusion >>
rect 43 -162 48 -156
rect 47 -166 48 -162
rect 50 -160 51 -156
rect 50 -166 55 -160
rect -27 -186 -26 -182
rect -31 -202 -26 -186
rect -24 -202 -16 -182
rect -14 -198 -9 -182
rect 3 -188 8 -182
rect 7 -192 8 -188
rect 10 -186 12 -182
rect 16 -186 18 -182
rect 10 -192 18 -186
rect 20 -188 25 -182
rect 20 -192 21 -188
rect 67 -188 72 -182
rect 71 -192 72 -188
rect 74 -186 76 -182
rect 80 -186 82 -182
rect 74 -192 82 -186
rect 84 -188 89 -182
rect 95 -184 100 -178
rect 99 -188 100 -184
rect 102 -182 103 -178
rect 102 -188 107 -182
rect 84 -192 85 -188
rect -14 -202 -13 -198
rect 116 -200 121 -184
rect 120 -204 121 -200
rect 123 -204 131 -184
rect 133 -188 134 -184
rect 133 -204 138 -188
rect -17 -247 -11 -243
rect -17 -248 -7 -247
rect 13 -247 16 -243
rect 6 -248 16 -247
rect -17 -251 -7 -250
rect -13 -255 -7 -251
rect 6 -251 16 -250
rect 6 -255 12 -251
rect -85 -268 -84 -264
rect -89 -274 -84 -268
rect -82 -268 -80 -264
rect -76 -268 -75 -264
rect -82 -274 -75 -268
rect -73 -270 -68 -264
rect -73 -274 -72 -270
rect 67 -270 72 -264
rect 71 -274 72 -270
rect 74 -268 75 -264
rect 79 -268 81 -264
rect 74 -274 81 -268
rect 83 -268 84 -264
rect 83 -274 88 -268
<< pdiffusion >>
rect 7 -128 8 -124
rect -27 -148 -26 -144
rect -31 -164 -26 -148
rect -24 -160 -16 -144
rect -24 -164 -22 -160
rect -18 -164 -16 -160
rect -14 -148 -13 -144
rect -14 -164 -9 -148
rect 3 -164 8 -128
rect 10 -164 18 -124
rect 20 -160 25 -124
rect 47 -128 48 -124
rect 43 -144 48 -128
rect 50 -140 55 -124
rect 50 -144 51 -140
rect 71 -128 72 -124
rect 20 -164 21 -160
rect 67 -164 72 -128
rect 74 -164 82 -124
rect 84 -160 89 -124
rect 84 -164 85 -160
rect 99 -150 100 -146
rect 95 -166 100 -150
rect 102 -162 107 -146
rect 102 -166 103 -162
rect 120 -150 121 -146
rect 116 -166 121 -150
rect 123 -162 131 -146
rect 123 -166 125 -162
rect 129 -166 131 -162
rect 133 -150 134 -146
rect 133 -166 138 -150
rect -89 -247 -84 -231
rect -85 -251 -84 -247
rect -82 -245 -75 -231
rect -82 -249 -80 -245
rect -76 -249 -75 -245
rect -82 -251 -75 -249
rect -73 -235 -72 -231
rect -73 -251 -68 -235
rect 71 -235 72 -231
rect -44 -247 -29 -242
rect -49 -248 -29 -247
rect 28 -247 43 -242
rect 28 -248 48 -247
rect -49 -251 -29 -250
rect -49 -255 -33 -251
rect 28 -251 48 -250
rect 67 -251 72 -235
rect 74 -245 81 -231
rect 74 -249 75 -245
rect 79 -249 81 -245
rect 74 -251 81 -249
rect 83 -247 88 -231
rect 83 -251 84 -247
rect 32 -255 48 -251
<< ndcontact >>
rect 43 -166 47 -162
rect 51 -160 55 -156
rect -31 -186 -27 -182
rect 3 -192 7 -188
rect 12 -186 16 -182
rect 21 -192 25 -188
rect 67 -192 71 -188
rect 76 -186 80 -182
rect 95 -188 99 -184
rect 103 -182 107 -178
rect 85 -192 89 -188
rect -13 -202 -9 -198
rect 116 -204 120 -200
rect 134 -188 138 -184
rect -11 -247 -7 -243
rect 6 -247 13 -243
rect -17 -255 -13 -251
rect 12 -255 16 -251
rect -89 -268 -85 -264
rect -80 -268 -76 -264
rect -72 -274 -68 -270
rect 67 -274 71 -270
rect 75 -268 79 -264
rect 84 -268 88 -264
<< pdcontact >>
rect 3 -128 7 -124
rect -31 -148 -27 -144
rect -22 -164 -18 -160
rect -13 -148 -9 -144
rect 43 -128 47 -124
rect 51 -144 55 -140
rect 67 -128 71 -124
rect 21 -164 25 -160
rect 85 -164 89 -160
rect 95 -150 99 -146
rect 103 -166 107 -162
rect 116 -150 120 -146
rect 125 -166 129 -162
rect 134 -150 138 -146
rect -89 -251 -85 -247
rect -80 -249 -76 -245
rect -72 -235 -68 -231
rect 67 -235 71 -231
rect -33 -255 -29 -251
rect 75 -249 79 -245
rect 84 -251 88 -247
rect 28 -255 32 -251
<< polysilicon >>
rect 8 -124 10 -121
rect 18 -124 20 -121
rect 48 -124 50 -120
rect 72 -124 74 -121
rect 82 -124 84 -121
rect -26 -144 -24 -140
rect -16 -144 -14 -140
rect 48 -156 50 -144
rect -26 -182 -24 -164
rect -16 -182 -14 -164
rect 8 -182 10 -164
rect 18 -182 20 -164
rect 100 -146 102 -143
rect 121 -146 123 -142
rect 131 -146 133 -142
rect 48 -170 50 -166
rect 72 -182 74 -164
rect 82 -182 84 -164
rect 100 -178 102 -166
rect 121 -184 123 -166
rect 131 -184 133 -166
rect 100 -191 102 -188
rect 8 -195 10 -192
rect 18 -195 20 -192
rect 72 -195 74 -192
rect 82 -195 84 -192
rect -26 -206 -24 -202
rect -16 -206 -14 -202
rect 121 -208 123 -204
rect 131 -208 133 -204
rect -84 -231 -82 -219
rect -75 -231 -73 -228
rect 72 -231 74 -228
rect 81 -231 83 -219
rect -53 -250 -49 -248
rect -29 -250 -17 -248
rect -7 -250 -3 -248
rect 2 -250 6 -248
rect 16 -250 28 -248
rect 48 -250 52 -248
rect -84 -257 -82 -251
rect -84 -264 -82 -260
rect -75 -264 -73 -251
rect 72 -264 74 -251
rect 81 -257 83 -251
rect 81 -264 83 -260
rect -84 -276 -82 -274
rect -84 -280 -83 -276
rect -75 -277 -73 -274
rect 72 -277 74 -274
rect 81 -276 83 -274
rect 82 -280 83 -276
rect -84 -281 -82 -280
rect 81 -281 83 -280
<< polycontact >>
rect 44 -155 48 -151
rect -24 -181 -20 -177
rect -14 -175 -10 -171
rect 4 -181 8 -177
rect 14 -175 18 -171
rect 68 -181 72 -177
rect 78 -175 82 -171
rect 96 -177 100 -173
rect 117 -177 121 -173
rect 127 -183 131 -179
rect -82 -224 -78 -220
rect 77 -224 81 -220
rect -22 -248 -18 -244
rect 17 -248 21 -244
rect -73 -262 -69 -258
rect 68 -262 72 -258
rect -83 -280 -79 -276
rect 78 -280 82 -276
<< metal1 >>
rect -6 -115 -3 -114
rect 2 -115 98 -114
rect -6 -117 98 -115
rect -6 -134 -3 -117
rect 3 -124 6 -117
rect 43 -124 46 -117
rect 67 -124 70 -117
rect -37 -137 -3 -134
rect 95 -136 98 -117
rect -31 -144 -27 -137
rect -12 -144 -9 -137
rect 95 -139 144 -136
rect 52 -151 55 -144
rect 95 -146 98 -139
rect 116 -146 119 -139
rect 134 -146 138 -139
rect 37 -154 44 -151
rect -22 -165 -19 -164
rect -31 -168 -19 -165
rect -31 -177 -28 -168
rect -10 -174 14 -171
rect 22 -173 25 -164
rect 22 -176 28 -173
rect -50 -180 -28 -177
rect -31 -182 -28 -180
rect -20 -181 4 -178
rect 22 -178 25 -176
rect 13 -181 25 -178
rect 37 -178 40 -154
rect 52 -154 63 -151
rect 52 -156 55 -154
rect 43 -171 46 -166
rect 60 -171 63 -154
rect 43 -174 56 -171
rect 60 -174 78 -171
rect 37 -181 49 -178
rect -5 -182 0 -181
rect 13 -182 16 -181
rect -38 -206 -35 -189
rect 3 -196 6 -192
rect 22 -195 25 -192
rect -50 -209 -35 -206
rect -12 -207 -9 -202
rect -6 -199 22 -196
rect -6 -207 -3 -199
rect -50 -221 -47 -209
rect -12 -210 -3 -207
rect -78 -224 -47 -221
rect -59 -231 -56 -224
rect -68 -234 -19 -231
rect -2 -234 1 -218
rect -88 -258 -85 -251
rect -22 -244 -19 -234
rect -4 -238 3 -234
rect 11 -243 14 -199
rect 46 -202 49 -181
rect 53 -194 56 -174
rect 86 -173 89 -164
rect 104 -173 107 -166
rect 126 -167 129 -166
rect 126 -170 138 -167
rect 86 -176 96 -173
rect 65 -180 68 -177
rect 86 -178 89 -176
rect 104 -176 117 -173
rect 104 -178 107 -176
rect 77 -181 89 -178
rect 77 -182 80 -181
rect 135 -179 138 -170
rect 115 -183 127 -180
rect 135 -182 144 -179
rect 135 -184 138 -182
rect 67 -196 70 -192
rect 86 -196 89 -192
rect 95 -195 98 -188
rect 57 -199 94 -196
rect 46 -205 61 -202
rect 58 -211 61 -205
rect 116 -208 119 -204
rect 120 -212 141 -209
rect 44 -223 45 -218
rect 50 -221 51 -218
rect 50 -223 77 -221
rect 44 -224 77 -223
rect 44 -225 51 -224
rect 55 -231 58 -224
rect -7 -246 6 -243
rect 13 -247 14 -243
rect 18 -234 67 -231
rect 18 -244 21 -234
rect -80 -252 -77 -249
rect -29 -255 -17 -252
rect 16 -255 28 -252
rect 76 -252 79 -249
rect -97 -260 -85 -258
rect -92 -261 -85 -260
rect -88 -264 -85 -261
rect -80 -264 -77 -257
rect -69 -262 -63 -259
rect -22 -263 -19 -255
rect -52 -266 -19 -263
rect 18 -263 21 -255
rect 62 -262 68 -259
rect 18 -266 51 -263
rect 76 -264 79 -257
rect -52 -269 -49 -266
rect -65 -271 -49 -269
rect -68 -272 -49 -271
rect 48 -269 51 -266
rect 84 -258 87 -251
rect 84 -260 96 -258
rect 84 -261 91 -260
rect 84 -264 87 -261
rect 48 -271 64 -269
rect 48 -272 67 -271
rect -68 -274 -62 -272
rect -65 -277 -62 -274
rect -79 -280 -62 -277
rect 61 -274 67 -272
rect 61 -277 64 -274
rect 61 -280 78 -277
<< m2contact >>
rect -46 -170 -40 -165
rect -55 -181 -50 -176
rect -5 -171 0 -166
rect 28 -177 33 -172
rect -39 -189 -34 -184
rect -5 -187 0 -182
rect -63 -216 -58 -211
rect -9 -239 -4 -234
rect 3 -239 8 -234
rect 22 -200 27 -195
rect 60 -182 65 -177
rect 110 -185 115 -180
rect 52 -199 57 -194
rect 94 -200 99 -195
rect 57 -216 62 -211
rect 115 -213 120 -208
rect -81 -257 -76 -252
rect 75 -257 80 -252
<< pdm12contact >>
rect -49 -247 -44 -242
rect 43 -247 48 -242
<< metal2 >>
rect -54 -160 114 -157
rect -54 -176 -51 -160
rect -40 -169 -5 -166
rect -46 -201 -43 -170
rect 29 -178 33 -177
rect 29 -181 60 -178
rect 111 -180 114 -160
rect -34 -187 -5 -184
rect 27 -199 52 -196
rect 99 -199 115 -196
rect -54 -204 -43 -201
rect -54 -212 -51 -204
rect -58 -215 -51 -212
rect -101 -253 -98 -225
rect -101 -256 -81 -253
rect -62 -258 -59 -216
rect 112 -212 115 -199
rect -48 -230 -13 -227
rect -48 -242 -45 -230
rect -16 -235 -13 -230
rect 12 -230 47 -227
rect -16 -238 -9 -235
rect 12 -235 15 -230
rect 8 -238 15 -235
rect 44 -242 47 -230
rect 58 -258 61 -216
rect 80 -256 103 -253
rect 100 -282 103 -256
<< m3contact >>
rect -102 -225 -97 -220
<< m123contact >>
rect -3 -115 2 -110
rect -3 -218 2 -213
rect 45 -223 50 -218
rect -97 -265 -92 -260
rect -63 -263 -58 -258
rect 57 -263 62 -258
rect 91 -265 96 -260
<< metal3 >>
rect -2 -213 1 -115
rect -103 -220 -96 -219
rect -103 -225 -102 -220
rect -97 -222 -96 -220
rect 44 -222 45 -218
rect -97 -223 45 -222
rect 50 -223 51 -218
rect -97 -225 51 -223
rect -103 -226 -96 -225
rect -95 -260 -63 -259
rect -92 -262 -63 -260
rect 62 -260 94 -259
rect 62 -262 91 -260
<< labels >>
rlabel metal1 -1 -236 -1 -236 3 vdd
rlabel metal1 -1 -244 -1 -244 3 gnd
rlabel metal1 -15 -136 -15 -136 5 vdd
rlabel metal1 14 -197 14 -197 1 gnd
rlabel metal1 4 -116 4 -115 5 vdd
rlabel metal1 138 -182 144 -179 7 c1
rlabel metal1 131 -211 131 -211 1 gnd
rlabel metal1 122 -138 122 -138 5 vdd
rlabel m2contact 61 -179 65 -178 1 p0_inv
rlabel metal1 105 -175 107 -172 1 temp100
rlabel metal1 68 -116 68 -115 5 vdd
rlabel metal1 78 -197 78 -197 1 gnd
rlabel metal1 53 -153 55 -150 1 c0_inv
rlabel metal1 38 -154 40 -152 3 c0
rlabel metal1 44 -173 44 -173 1 gnd
rlabel metal1 43 -115 43 -115 5 vdd
rlabel m2contact 59 -214 60 -214 1 c0
rlabel metal2 101 -282 102 -280 1 s0
rlabel metal2 -100 -255 -96 -253 3 mid_s0
rlabel metal1 -8 -174 3 -171 1 a0
rlabel metal1 -8 -181 3 -178 1 b0
rlabel metal1 -37 -180 -31 -177 1 g0_inv
rlabel metal1 25 -176 30 -173 1 p0_inv
rlabel m2contact 111 -183 115 -181 1 g0_inv
<< end >>
