* SPICE3 file created from NOR.ext - technology: scmos
* NOR gate layout
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global gnd vdd

M1000 out in2 a_n11_40# w_n24_34# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1001 out in1 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=100 ps=60
M1002 a_n11_40# in1 vdd w_n24_34# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1003 gnd in2 out Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in1 in2 0.24fF
C1 w_n24_34# vdd 0.02fF
C2 out gnd 0.02fF
C3 w_n24_34# out 0.02fF
C4 w_n24_34# in2 0.06fF
C5 in2 out 0.17fF
C6 in1 gnd 0.02fF
C7 w_n24_34# in1 0.06fF
C8 in1 out 0.02fF
C9 gnd Gnd 0.10fF
C10 out Gnd 0.07fF
C11 vdd Gnd 0.09fF
C12 in2 Gnd 0.18fF
C13 in1 Gnd 0.16fF
C14 w_n24_34# Gnd 1.78fF

Vdd vdd gnd 'SUPPLY'
Vin1 in1 gnd pulse 0 1.8 0 0.01ns 0.01ns 10ns 20ns
Vin2 in2 gnd pulse 0 1.8 0 0.01ns 0.01ns 20ns 40ns

.tran 1p 50n

.control
set hcopypscolor = 1
set color0=white
set color1=black

run

set curplottitle="2023112005_NOR"
plot v(in1), v(in2)+2, v(out)+4
.endc