magic
tech scmos
timestamp 1731382288
<< nwell >>
rect -158 94 -134 126
rect -110 94 -86 126
rect -63 100 -15 132
<< ntransistor >>
rect -147 66 -145 86
rect -123 59 -121 79
rect -99 66 -97 86
rect -75 59 -73 79
rect -52 69 -50 89
rect -28 69 -26 89
<< ptransistor >>
rect -147 100 -145 120
rect -99 100 -97 120
rect -52 106 -50 126
rect -28 106 -26 126
<< ndiffusion >>
rect -152 70 -147 86
rect -148 66 -147 70
rect -145 70 -140 86
rect -145 66 -144 70
rect -124 75 -123 79
rect -128 59 -123 75
rect -121 63 -116 79
rect -104 70 -99 86
rect -100 66 -99 70
rect -97 70 -92 86
rect -97 66 -96 70
rect -76 75 -75 79
rect -121 59 -120 63
rect -80 59 -75 75
rect -73 63 -68 79
rect -57 73 -52 89
rect -53 69 -52 73
rect -50 85 -49 89
rect -50 69 -45 85
rect -33 73 -28 89
rect -29 69 -28 73
rect -26 85 -25 89
rect -26 69 -21 85
rect -73 59 -72 63
<< pdiffusion >>
rect -53 122 -52 126
rect -148 116 -147 120
rect -152 100 -147 116
rect -145 104 -140 120
rect -145 100 -144 104
rect -100 116 -99 120
rect -104 100 -99 116
rect -97 104 -92 120
rect -57 106 -52 122
rect -50 110 -45 126
rect -50 106 -49 110
rect -29 122 -28 126
rect -33 106 -28 122
rect -26 110 -21 126
rect -26 106 -25 110
rect -97 100 -96 104
<< ndcontact >>
rect -152 66 -148 70
rect -144 66 -140 70
rect -128 75 -124 79
rect -104 66 -100 70
rect -96 66 -92 70
rect -80 75 -76 79
rect -120 59 -116 63
rect -57 69 -53 73
rect -49 85 -45 89
rect -33 69 -29 73
rect -25 85 -21 89
rect -72 59 -68 63
<< pdcontact >>
rect -57 122 -53 126
rect -152 116 -148 120
rect -144 100 -140 104
rect -104 116 -100 120
rect -49 106 -45 110
rect -33 122 -29 126
rect -25 106 -21 110
rect -96 100 -92 104
<< polysilicon >>
rect -52 126 -50 129
rect -28 126 -26 129
rect -147 120 -145 123
rect -99 120 -97 123
rect -147 86 -145 100
rect -123 79 -121 91
rect -99 86 -97 100
rect -147 62 -145 66
rect -75 79 -73 91
rect -52 89 -50 106
rect -28 89 -26 106
rect -99 62 -97 66
rect -52 65 -50 69
rect -28 65 -26 69
rect -123 56 -121 59
rect -75 56 -73 59
<< polycontact >>
rect -151 89 -147 93
rect -127 85 -123 89
rect -103 89 -99 93
rect -56 93 -52 97
rect -79 85 -75 89
rect -32 93 -28 97
<< metal1 >>
rect -97 135 -19 138
rect -97 131 -94 135
rect -158 128 -94 131
rect -152 120 -149 128
rect -104 120 -101 128
rect -57 126 -54 135
rect -33 126 -30 135
rect -160 89 -151 92
rect -143 90 -140 100
rect -137 94 -112 97
rect -137 90 -134 94
rect -143 87 -134 90
rect -115 92 -112 94
rect -115 89 -103 92
rect -95 90 -92 100
rect -49 97 -45 106
rect -89 94 -56 97
rect -89 90 -86 94
rect -49 93 -32 97
rect -25 96 -21 106
rect -25 93 -15 96
rect -138 82 -134 87
rect -131 85 -127 88
rect -95 87 -86 90
rect -49 89 -45 93
rect -90 82 -86 87
rect -83 85 -79 88
rect -25 89 -21 93
rect -138 79 -125 82
rect -90 79 -77 82
rect -152 50 -149 66
rect -143 56 -140 66
rect -120 56 -117 59
rect -143 53 -117 56
rect -104 50 -101 66
rect -95 57 -92 66
rect -57 64 -54 69
rect -33 64 -30 69
rect -57 61 -30 64
rect -72 57 -69 59
rect -95 54 -69 57
rect -57 50 -54 61
rect -152 47 -54 50
<< labels >>
rlabel metal1 -151 129 -151 129 5 vdd
rlabel metal1 -51 137 -50 137 5 vdd
rlabel metal1 -27 137 -26 137 5 vdd
rlabel metal1 -129 86 -129 86 1 clk
rlabel metal1 -157 91 -157 91 1 d
rlabel metal1 -81 86 -81 86 1 clk
rlabel metal1 -78 96 -77 96 1 q
rlabel metal1 -60 95 -60 95 3 in
rlabel metal1 -20 94 -20 94 7 out
rlabel metal1 -102 48 -102 48 1 gnd
<< end >>
