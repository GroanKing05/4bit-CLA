* SPICE3 file created from OR.ext - technology: scmos

.option scale=0.09u

M1000 out a_n11_12# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=150 ps=90
M1001 a_n11_12# in2 a_n11_40# w_n24_34# pfet w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1002 a_n11_12# in1 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1003 out a_n11_12# vdd w_n24_34# pfet w=20 l=2
+  ad=100 pd=50 as=300 ps=140
M1004 a_n11_40# in1 vdd w_n24_34# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 gnd in2 a_n11_12# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n24_34# in2 0.06fF
C1 in2 a_n11_12# 0.17fF
C2 w_n24_34# in1 0.06fF
C3 a_n11_12# gnd 0.04fF
C4 in1 a_n11_12# 0.02fF
C5 w_n24_34# out 0.02fF
C6 w_n24_34# vdd 0.07fF
C7 in1 in2 0.24fF
C8 a_n11_12# out 0.04fF
C9 in1 gnd 0.02fF
C10 w_n24_34# a_n11_12# 0.09fF
C11 gnd Gnd 0.14fF
C12 out Gnd 0.03fF
C13 a_n11_12# Gnd 0.18fF
C14 vdd Gnd 0.17fF
C15 in2 Gnd 0.18fF
C16 in1 Gnd 0.16fF
C17 w_n24_34# Gnd 2.40fF
