magic
tech scmos
timestamp 1731411278
<< nwell >>
rect 293 -83 325 -64
rect 293 -89 347 -83
rect 295 -117 347 -89
rect 365 -99 442 -77
rect 365 -109 460 -99
rect -3 -138 31 -118
rect -37 -170 31 -138
rect 37 -140 95 -118
rect 37 -150 144 -140
rect 210 -144 244 -124
rect 272 -137 306 -131
rect 61 -170 144 -150
rect 89 -172 144 -170
rect 176 -176 244 -144
rect 250 -163 306 -137
rect 250 -169 275 -163
rect 323 -177 357 -125
rect 408 -129 460 -109
rect 436 -131 460 -129
rect -95 -257 -62 -225
rect -55 -262 -23 -236
rect 22 -262 54 -236
rect 61 -257 94 -225
rect 118 -263 151 -231
rect 158 -268 190 -242
rect 235 -268 267 -242
rect 274 -263 307 -231
<< ntransistor >>
rect 277 -78 287 -76
rect 273 -96 283 -94
rect 273 -106 283 -104
rect 48 -166 50 -156
rect -26 -202 -24 -182
rect -16 -202 -14 -182
rect 8 -192 10 -182
rect 18 -192 20 -182
rect 72 -192 74 -182
rect 82 -192 84 -182
rect 100 -188 102 -178
rect 121 -204 123 -184
rect 131 -204 133 -184
rect 376 -141 378 -121
rect 386 -141 388 -121
rect 419 -151 421 -141
rect 429 -151 431 -141
rect 447 -147 449 -137
rect 262 -185 264 -175
rect 187 -208 189 -188
rect 197 -208 199 -188
rect 221 -198 223 -188
rect 231 -198 233 -188
rect 283 -195 285 -175
rect 293 -195 295 -175
rect 334 -199 336 -189
rect 344 -199 346 -189
rect -17 -250 -7 -248
rect 6 -250 16 -248
rect 196 -256 206 -254
rect 219 -256 229 -254
rect -84 -274 -82 -264
rect -75 -274 -73 -264
rect 72 -274 74 -264
rect 81 -274 83 -264
rect 129 -280 131 -270
rect 138 -280 140 -270
rect 285 -280 287 -270
rect 294 -280 296 -270
<< ptransistor >>
rect 299 -78 319 -76
rect 301 -96 341 -94
rect 376 -103 378 -83
rect 386 -103 388 -83
rect 301 -106 341 -104
rect -26 -164 -24 -144
rect -16 -164 -14 -144
rect 8 -164 10 -124
rect 18 -164 20 -124
rect 48 -144 50 -124
rect 72 -164 74 -124
rect 82 -164 84 -124
rect 100 -166 102 -146
rect 121 -166 123 -146
rect 131 -166 133 -146
rect 187 -170 189 -150
rect 197 -170 199 -150
rect 221 -170 223 -130
rect 231 -170 233 -130
rect 262 -163 264 -143
rect 283 -157 285 -137
rect 293 -157 295 -137
rect 334 -171 336 -131
rect 344 -171 346 -131
rect 419 -123 421 -83
rect 429 -123 431 -83
rect 447 -125 449 -105
rect -84 -251 -82 -231
rect -75 -251 -73 -231
rect -49 -250 -29 -248
rect 28 -250 48 -248
rect 72 -251 74 -231
rect 81 -251 83 -231
rect 129 -257 131 -237
rect 138 -257 140 -237
rect 164 -256 184 -254
rect 241 -256 261 -254
rect 285 -257 287 -237
rect 294 -257 296 -237
<< ndiffusion >>
rect 277 -75 283 -71
rect 277 -76 287 -75
rect 277 -79 287 -78
rect 281 -83 287 -79
rect 277 -93 283 -89
rect 273 -94 283 -93
rect 273 -98 283 -96
rect 273 -102 279 -98
rect 273 -104 283 -102
rect 273 -107 283 -106
rect 277 -111 283 -107
rect 43 -162 48 -156
rect 47 -166 48 -162
rect 50 -160 51 -156
rect 50 -166 55 -160
rect -27 -186 -26 -182
rect -31 -202 -26 -186
rect -24 -202 -16 -182
rect -14 -198 -9 -182
rect 3 -188 8 -182
rect 7 -192 8 -188
rect 10 -186 12 -182
rect 16 -186 18 -182
rect 10 -192 18 -186
rect 20 -188 25 -182
rect 20 -192 21 -188
rect 67 -188 72 -182
rect 71 -192 72 -188
rect 74 -186 76 -182
rect 80 -186 82 -182
rect 74 -192 82 -186
rect 84 -188 89 -182
rect 95 -184 100 -178
rect 99 -188 100 -184
rect 102 -182 103 -178
rect 102 -188 107 -182
rect 84 -192 85 -188
rect -14 -202 -13 -198
rect 116 -200 121 -184
rect 120 -204 121 -200
rect 123 -204 131 -184
rect 133 -188 134 -184
rect 371 -137 376 -121
rect 375 -141 376 -137
rect 378 -141 386 -121
rect 388 -125 389 -121
rect 388 -141 393 -125
rect 414 -147 419 -141
rect 418 -151 419 -147
rect 421 -145 423 -141
rect 427 -145 429 -141
rect 421 -151 429 -145
rect 431 -147 436 -141
rect 442 -143 447 -137
rect 446 -147 447 -143
rect 449 -141 450 -137
rect 449 -147 454 -141
rect 431 -151 432 -147
rect 261 -179 262 -175
rect 257 -185 262 -179
rect 264 -181 269 -175
rect 264 -185 265 -181
rect 282 -179 283 -175
rect 133 -204 138 -188
rect 186 -192 187 -188
rect 182 -208 187 -192
rect 189 -208 197 -188
rect 199 -204 204 -188
rect 216 -194 221 -188
rect 220 -198 221 -194
rect 223 -192 225 -188
rect 229 -192 231 -188
rect 223 -198 231 -192
rect 233 -194 238 -188
rect 233 -198 234 -194
rect 278 -195 283 -179
rect 285 -195 293 -175
rect 295 -191 300 -175
rect 295 -195 296 -191
rect 329 -195 334 -189
rect 333 -199 334 -195
rect 336 -193 338 -189
rect 342 -193 344 -189
rect 336 -199 344 -193
rect 346 -195 351 -189
rect 346 -199 347 -195
rect 199 -208 200 -204
rect -17 -247 -11 -243
rect -17 -248 -7 -247
rect 13 -247 16 -243
rect 6 -248 16 -247
rect -17 -251 -7 -250
rect -13 -255 -7 -251
rect 6 -251 16 -250
rect 6 -255 12 -251
rect 196 -253 202 -249
rect 196 -254 206 -253
rect 226 -253 229 -249
rect 219 -254 229 -253
rect -85 -268 -84 -264
rect -89 -274 -84 -268
rect -82 -268 -80 -264
rect -76 -268 -75 -264
rect -82 -274 -75 -268
rect -73 -270 -68 -264
rect -73 -274 -72 -270
rect 67 -270 72 -264
rect 71 -274 72 -270
rect 74 -268 75 -264
rect 79 -268 81 -264
rect 74 -274 81 -268
rect 83 -268 84 -264
rect 83 -274 88 -268
rect 196 -257 206 -256
rect 200 -261 206 -257
rect 219 -257 229 -256
rect 219 -261 225 -257
rect 128 -274 129 -270
rect 124 -280 129 -274
rect 131 -274 133 -270
rect 137 -274 138 -270
rect 131 -280 138 -274
rect 140 -276 145 -270
rect 140 -280 141 -276
rect 280 -276 285 -270
rect 284 -280 285 -276
rect 287 -274 288 -270
rect 292 -274 294 -270
rect 287 -280 294 -274
rect 296 -274 297 -270
rect 296 -280 301 -274
<< pdiffusion >>
rect 303 -75 319 -71
rect 299 -76 319 -75
rect 299 -79 319 -78
rect 299 -83 315 -79
rect 375 -87 376 -83
rect 305 -93 341 -89
rect 301 -94 341 -93
rect 301 -104 341 -96
rect 371 -103 376 -87
rect 378 -99 386 -83
rect 378 -103 380 -99
rect 384 -103 386 -99
rect 388 -87 389 -83
rect 388 -103 393 -87
rect 418 -87 419 -83
rect 301 -107 341 -106
rect 301 -111 337 -107
rect 7 -128 8 -124
rect -27 -148 -26 -144
rect -31 -164 -26 -148
rect -24 -160 -16 -144
rect -24 -164 -22 -160
rect -18 -164 -16 -160
rect -14 -148 -13 -144
rect -14 -164 -9 -148
rect 3 -164 8 -128
rect 10 -164 18 -124
rect 20 -160 25 -124
rect 47 -128 48 -124
rect 43 -144 48 -128
rect 50 -140 55 -124
rect 50 -144 51 -140
rect 71 -128 72 -124
rect 20 -164 21 -160
rect 67 -164 72 -128
rect 74 -164 82 -124
rect 84 -160 89 -124
rect 220 -134 221 -130
rect 84 -164 85 -160
rect 99 -150 100 -146
rect 95 -166 100 -150
rect 102 -162 107 -146
rect 102 -166 103 -162
rect 120 -150 121 -146
rect 116 -166 121 -150
rect 123 -162 131 -146
rect 123 -166 125 -162
rect 129 -166 131 -162
rect 133 -150 134 -146
rect 133 -166 138 -150
rect 186 -154 187 -150
rect 182 -170 187 -154
rect 189 -166 197 -150
rect 189 -170 191 -166
rect 195 -170 197 -166
rect 199 -154 200 -150
rect 199 -170 204 -154
rect 216 -170 221 -134
rect 223 -170 231 -130
rect 233 -166 238 -130
rect 282 -141 283 -137
rect 257 -159 262 -143
rect 261 -163 262 -159
rect 264 -147 265 -143
rect 264 -163 269 -147
rect 278 -157 283 -141
rect 285 -153 293 -137
rect 285 -157 287 -153
rect 291 -157 293 -153
rect 295 -141 296 -137
rect 295 -157 300 -141
rect 233 -170 234 -166
rect 329 -167 334 -131
rect 333 -171 334 -167
rect 336 -171 344 -131
rect 346 -135 347 -131
rect 346 -171 351 -135
rect 414 -123 419 -87
rect 421 -123 429 -83
rect 431 -119 436 -83
rect 431 -123 432 -119
rect 446 -109 447 -105
rect 442 -125 447 -109
rect 449 -121 454 -105
rect 449 -125 450 -121
rect -89 -247 -84 -231
rect -85 -251 -84 -247
rect -82 -245 -75 -231
rect -82 -249 -80 -245
rect -76 -249 -75 -245
rect -82 -251 -75 -249
rect -73 -235 -72 -231
rect -73 -251 -68 -235
rect 71 -235 72 -231
rect -44 -247 -29 -242
rect -49 -248 -29 -247
rect 28 -247 43 -242
rect 28 -248 48 -247
rect -49 -251 -29 -250
rect -49 -255 -33 -251
rect 28 -251 48 -250
rect 67 -251 72 -235
rect 74 -245 81 -231
rect 74 -249 75 -245
rect 79 -249 81 -245
rect 74 -251 81 -249
rect 83 -247 88 -231
rect 83 -251 84 -247
rect 32 -255 48 -251
rect 124 -253 129 -237
rect 128 -257 129 -253
rect 131 -251 138 -237
rect 131 -255 133 -251
rect 137 -255 138 -251
rect 131 -257 138 -255
rect 140 -241 141 -237
rect 140 -257 145 -241
rect 284 -241 285 -237
rect 169 -253 184 -248
rect 164 -254 184 -253
rect 241 -253 256 -248
rect 241 -254 261 -253
rect 164 -257 184 -256
rect 164 -261 180 -257
rect 241 -257 261 -256
rect 280 -257 285 -241
rect 287 -251 294 -237
rect 287 -255 288 -251
rect 292 -255 294 -251
rect 287 -257 294 -255
rect 296 -253 301 -237
rect 296 -257 297 -253
rect 245 -261 261 -257
<< ndcontact >>
rect 283 -75 287 -71
rect 277 -83 281 -79
rect 273 -93 277 -89
rect 279 -102 283 -98
rect 273 -111 277 -107
rect 43 -166 47 -162
rect 51 -160 55 -156
rect -31 -186 -27 -182
rect 3 -192 7 -188
rect 12 -186 16 -182
rect 21 -192 25 -188
rect 67 -192 71 -188
rect 76 -186 80 -182
rect 95 -188 99 -184
rect 103 -182 107 -178
rect 85 -192 89 -188
rect -13 -202 -9 -198
rect 116 -204 120 -200
rect 134 -188 138 -184
rect 371 -141 375 -137
rect 389 -125 393 -121
rect 414 -151 418 -147
rect 423 -145 427 -141
rect 442 -147 446 -143
rect 450 -141 454 -137
rect 432 -151 436 -147
rect 257 -179 261 -175
rect 265 -185 269 -181
rect 278 -179 282 -175
rect 182 -192 186 -188
rect 216 -198 220 -194
rect 225 -192 229 -188
rect 234 -198 238 -194
rect 296 -195 300 -191
rect 329 -199 333 -195
rect 338 -193 342 -189
rect 347 -199 351 -195
rect 200 -208 204 -204
rect -11 -247 -7 -243
rect 6 -247 13 -243
rect -17 -255 -13 -251
rect 12 -255 16 -251
rect 202 -253 206 -249
rect 219 -253 226 -249
rect -89 -268 -85 -264
rect -80 -268 -76 -264
rect -72 -274 -68 -270
rect 67 -274 71 -270
rect 75 -268 79 -264
rect 84 -268 88 -264
rect 196 -261 200 -257
rect 225 -261 229 -257
rect 124 -274 128 -270
rect 133 -274 137 -270
rect 141 -280 145 -276
rect 280 -280 284 -276
rect 288 -274 292 -270
rect 297 -274 301 -270
<< pdcontact >>
rect 299 -75 303 -71
rect 315 -83 319 -79
rect 371 -87 375 -83
rect 301 -93 305 -89
rect 380 -103 384 -99
rect 389 -87 393 -83
rect 414 -87 418 -83
rect 337 -111 341 -107
rect 3 -128 7 -124
rect -31 -148 -27 -144
rect -22 -164 -18 -160
rect -13 -148 -9 -144
rect 43 -128 47 -124
rect 51 -144 55 -140
rect 67 -128 71 -124
rect 21 -164 25 -160
rect 216 -134 220 -130
rect 85 -164 89 -160
rect 95 -150 99 -146
rect 103 -166 107 -162
rect 116 -150 120 -146
rect 125 -166 129 -162
rect 134 -150 138 -146
rect 182 -154 186 -150
rect 191 -170 195 -166
rect 200 -154 204 -150
rect 278 -141 282 -137
rect 257 -163 261 -159
rect 265 -147 269 -143
rect 287 -157 291 -153
rect 296 -141 300 -137
rect 234 -170 238 -166
rect 329 -171 333 -167
rect 347 -135 351 -131
rect 432 -123 436 -119
rect 442 -109 446 -105
rect 450 -125 454 -121
rect -89 -251 -85 -247
rect -80 -249 -76 -245
rect -72 -235 -68 -231
rect 67 -235 71 -231
rect -33 -255 -29 -251
rect 75 -249 79 -245
rect 84 -251 88 -247
rect 28 -255 32 -251
rect 124 -257 128 -253
rect 133 -255 137 -251
rect 141 -241 145 -237
rect 280 -241 284 -237
rect 180 -261 184 -257
rect 288 -255 292 -251
rect 297 -257 301 -253
rect 241 -261 245 -257
<< polysilicon >>
rect 274 -78 277 -76
rect 287 -78 299 -76
rect 319 -78 322 -76
rect 376 -83 378 -79
rect 386 -83 388 -79
rect 419 -83 421 -80
rect 429 -83 431 -80
rect 270 -96 273 -94
rect 283 -96 301 -94
rect 341 -96 344 -94
rect 270 -106 273 -104
rect 283 -106 301 -104
rect 341 -106 344 -104
rect 8 -124 10 -121
rect 18 -124 20 -121
rect 48 -124 50 -120
rect 376 -121 378 -103
rect 386 -121 388 -103
rect 72 -124 74 -121
rect 82 -124 84 -121
rect -26 -144 -24 -140
rect -16 -144 -14 -140
rect 48 -156 50 -144
rect -26 -182 -24 -164
rect -16 -182 -14 -164
rect 8 -182 10 -164
rect 18 -182 20 -164
rect 221 -130 223 -127
rect 231 -130 233 -127
rect 100 -146 102 -143
rect 121 -146 123 -142
rect 131 -146 133 -142
rect 48 -170 50 -166
rect 72 -182 74 -164
rect 82 -182 84 -164
rect 187 -150 189 -146
rect 197 -150 199 -146
rect 100 -178 102 -166
rect 121 -184 123 -166
rect 131 -184 133 -166
rect 334 -131 336 -128
rect 344 -131 346 -128
rect 283 -137 285 -133
rect 293 -137 295 -133
rect 262 -143 264 -139
rect 100 -191 102 -188
rect 8 -195 10 -192
rect 18 -195 20 -192
rect 72 -195 74 -192
rect 82 -195 84 -192
rect -26 -206 -24 -202
rect -16 -206 -14 -202
rect 187 -188 189 -170
rect 197 -188 199 -170
rect 221 -188 223 -170
rect 231 -188 233 -170
rect 262 -175 264 -163
rect 283 -175 285 -157
rect 293 -175 295 -157
rect 447 -105 449 -102
rect 419 -141 421 -123
rect 429 -141 431 -123
rect 447 -137 449 -125
rect 376 -145 378 -141
rect 386 -145 388 -141
rect 447 -150 449 -147
rect 419 -154 421 -151
rect 429 -154 431 -151
rect 121 -208 123 -204
rect 131 -208 133 -204
rect 262 -189 264 -185
rect 334 -189 336 -171
rect 344 -189 346 -171
rect 221 -201 223 -198
rect 231 -201 233 -198
rect 283 -199 285 -195
rect 293 -199 295 -195
rect 334 -202 336 -199
rect 344 -202 346 -199
rect 187 -212 189 -208
rect 197 -212 199 -208
rect -84 -231 -82 -219
rect -75 -231 -73 -228
rect 72 -231 74 -228
rect 81 -231 83 -219
rect -53 -250 -49 -248
rect -29 -250 -17 -248
rect -7 -250 -3 -248
rect 2 -250 6 -248
rect 16 -250 28 -248
rect 48 -250 52 -248
rect -84 -257 -82 -251
rect -84 -264 -82 -260
rect -75 -264 -73 -251
rect 129 -237 131 -225
rect 138 -237 140 -234
rect 285 -237 287 -234
rect 294 -237 296 -225
rect 72 -264 74 -251
rect 81 -257 83 -251
rect 160 -256 164 -254
rect 184 -256 196 -254
rect 206 -256 210 -254
rect 215 -256 219 -254
rect 229 -256 241 -254
rect 261 -256 265 -254
rect 81 -264 83 -260
rect 129 -263 131 -257
rect 129 -270 131 -266
rect 138 -270 140 -257
rect 285 -270 287 -257
rect 294 -263 296 -257
rect 294 -270 296 -266
rect -84 -276 -82 -274
rect -84 -280 -83 -276
rect -75 -277 -73 -274
rect 72 -277 74 -274
rect 81 -276 83 -274
rect 82 -280 83 -276
rect -84 -281 -82 -280
rect 81 -281 83 -280
rect 129 -282 131 -280
rect 129 -286 130 -282
rect 138 -283 140 -280
rect 285 -283 287 -280
rect 294 -282 296 -280
rect 295 -286 296 -282
rect 129 -287 131 -286
rect 294 -287 296 -286
<< polycontact >>
rect 288 -82 292 -78
rect 290 -100 294 -96
rect 284 -110 288 -106
rect 372 -114 376 -110
rect 382 -120 386 -116
rect 44 -155 48 -151
rect -24 -181 -20 -177
rect -14 -175 -10 -171
rect 4 -181 8 -177
rect 14 -175 18 -171
rect 68 -181 72 -177
rect 78 -175 82 -171
rect 96 -177 100 -173
rect 117 -177 121 -173
rect 127 -183 131 -179
rect 189 -187 193 -183
rect 199 -181 203 -177
rect 217 -187 221 -183
rect 227 -181 231 -177
rect 264 -174 268 -170
rect 285 -174 289 -170
rect 295 -168 299 -164
rect 415 -140 419 -136
rect 425 -134 429 -130
rect 443 -136 447 -132
rect 336 -182 340 -178
rect 346 -188 350 -184
rect -82 -224 -78 -220
rect 77 -224 81 -220
rect -22 -248 -18 -244
rect 17 -248 21 -244
rect 131 -230 135 -226
rect 290 -230 294 -226
rect -73 -262 -69 -258
rect 68 -262 72 -258
rect 191 -254 195 -250
rect 230 -254 234 -250
rect 140 -268 144 -264
rect 281 -268 285 -264
rect -83 -280 -79 -276
rect 78 -280 82 -276
rect 130 -286 134 -282
rect 291 -286 295 -282
<< metal1 >>
rect 289 -67 329 -64
rect 289 -71 292 -67
rect 287 -74 299 -71
rect 326 -73 329 -67
rect 326 -76 357 -73
rect 370 -76 445 -73
rect 266 -83 277 -80
rect 266 -89 269 -83
rect 289 -89 292 -82
rect 319 -83 346 -80
rect 266 -92 273 -89
rect 266 -107 269 -92
rect 284 -92 301 -89
rect 284 -98 287 -92
rect 283 -101 287 -98
rect -6 -115 -3 -114
rect 269 -111 273 -108
rect 2 -115 98 -114
rect 284 -115 288 -110
rect -6 -117 98 -115
rect -6 -134 -3 -117
rect 3 -124 6 -117
rect 43 -124 46 -117
rect 67 -124 70 -117
rect -37 -137 -3 -134
rect 95 -136 98 -117
rect 207 -121 210 -120
rect 291 -117 294 -100
rect 348 -108 351 -85
rect 341 -111 351 -108
rect 215 -121 272 -120
rect 207 -123 272 -121
rect 348 -121 351 -111
rect 354 -110 357 -76
rect 371 -83 374 -76
rect 389 -83 393 -76
rect 414 -83 417 -76
rect 381 -104 384 -103
rect 381 -107 393 -104
rect 354 -113 372 -110
rect 390 -116 393 -107
rect 442 -105 445 -76
rect 369 -120 382 -117
rect 390 -119 411 -116
rect 390 -121 393 -119
rect -31 -144 -27 -137
rect -12 -144 -9 -137
rect 95 -139 144 -136
rect 52 -151 55 -144
rect 95 -146 98 -139
rect 116 -146 119 -139
rect 134 -146 138 -139
rect 207 -140 210 -123
rect 216 -130 219 -123
rect 269 -127 272 -123
rect 303 -124 351 -121
rect 303 -127 306 -124
rect 266 -130 306 -127
rect 176 -143 210 -140
rect 266 -143 269 -130
rect 278 -137 282 -130
rect 297 -137 300 -130
rect 348 -131 351 -124
rect 408 -130 411 -119
rect 408 -133 425 -130
rect 433 -132 436 -123
rect 451 -132 454 -125
rect 433 -135 443 -132
rect 411 -139 415 -136
rect 433 -137 436 -135
rect 451 -135 461 -132
rect 451 -137 454 -135
rect 424 -140 436 -137
rect 424 -141 427 -140
rect 182 -150 186 -143
rect 201 -150 204 -143
rect 371 -146 374 -141
rect 37 -154 44 -151
rect -22 -165 -19 -164
rect -31 -168 -19 -165
rect -31 -177 -28 -168
rect -10 -174 14 -171
rect 22 -173 25 -164
rect 22 -176 28 -173
rect -50 -180 -28 -177
rect -31 -182 -28 -180
rect -20 -181 4 -178
rect 22 -178 25 -176
rect 13 -181 25 -178
rect 37 -178 40 -154
rect 52 -154 63 -151
rect 362 -149 410 -146
rect 52 -156 55 -154
rect 43 -171 46 -166
rect 60 -171 63 -154
rect 287 -158 290 -157
rect 43 -174 56 -171
rect 60 -174 78 -171
rect 37 -181 49 -178
rect -5 -182 0 -181
rect 13 -182 16 -181
rect -38 -206 -35 -189
rect 3 -196 6 -192
rect 22 -195 25 -192
rect -50 -209 -35 -206
rect -12 -207 -9 -202
rect -6 -199 22 -196
rect -6 -207 -3 -199
rect -50 -221 -47 -209
rect -12 -210 -3 -207
rect -78 -224 -47 -221
rect -59 -231 -56 -224
rect -68 -234 -19 -231
rect -2 -234 1 -218
rect -88 -258 -85 -251
rect -22 -244 -19 -234
rect -4 -238 3 -234
rect 11 -243 14 -199
rect 46 -202 49 -181
rect 53 -194 56 -174
rect 86 -173 89 -164
rect 278 -161 290 -158
rect 104 -173 107 -166
rect 126 -167 129 -166
rect 126 -170 138 -167
rect 86 -176 96 -173
rect 65 -180 68 -177
rect 86 -178 89 -176
rect 104 -176 117 -173
rect 104 -178 107 -176
rect 77 -181 89 -178
rect 77 -182 80 -181
rect 135 -179 138 -170
rect 257 -170 260 -163
rect 278 -170 281 -161
rect 299 -167 326 -164
rect 191 -171 194 -170
rect 182 -174 194 -171
rect 115 -183 127 -180
rect 135 -182 144 -179
rect 135 -184 138 -182
rect 67 -196 70 -192
rect 86 -196 89 -192
rect 95 -195 98 -188
rect 57 -199 94 -196
rect 141 -200 144 -182
rect 46 -205 61 -202
rect 58 -211 61 -205
rect 141 -203 157 -200
rect 116 -208 119 -204
rect 168 -206 171 -176
rect 182 -183 185 -174
rect 203 -180 227 -177
rect 235 -179 238 -170
rect 254 -173 260 -170
rect 257 -175 260 -173
rect 268 -173 281 -170
rect 278 -175 281 -173
rect 289 -174 308 -171
rect 235 -182 247 -179
rect 323 -180 326 -167
rect 329 -180 332 -171
rect 179 -186 185 -183
rect 182 -188 185 -186
rect 193 -187 217 -184
rect 235 -184 238 -182
rect 226 -187 238 -184
rect 244 -185 247 -182
rect 323 -183 332 -180
rect 340 -181 353 -178
rect 208 -188 213 -187
rect 226 -188 229 -187
rect 151 -209 171 -206
rect 120 -212 141 -209
rect 151 -217 154 -209
rect 175 -212 178 -195
rect 216 -202 219 -198
rect 235 -200 238 -198
rect 266 -199 269 -185
rect 329 -185 332 -183
rect 329 -188 341 -185
rect 350 -187 358 -184
rect 338 -189 341 -188
rect 235 -202 265 -200
rect 207 -203 265 -202
rect 163 -215 178 -212
rect 201 -213 204 -208
rect 207 -205 238 -203
rect 297 -200 300 -195
rect 270 -203 306 -200
rect 329 -203 332 -199
rect 348 -203 351 -199
rect 362 -203 365 -149
rect 407 -155 410 -149
rect 414 -155 417 -151
rect 433 -155 436 -151
rect 442 -155 445 -147
rect 407 -158 445 -155
rect 207 -213 210 -205
rect 44 -223 45 -218
rect 50 -221 51 -218
rect 50 -223 77 -221
rect 44 -224 77 -223
rect 44 -225 51 -224
rect 55 -231 58 -224
rect 163 -227 166 -215
rect 201 -216 210 -213
rect 135 -230 166 -227
rect -7 -246 6 -243
rect 13 -247 14 -243
rect 18 -234 67 -231
rect 18 -244 21 -234
rect 154 -237 157 -230
rect 145 -240 194 -237
rect 211 -240 214 -224
rect -80 -252 -77 -249
rect -29 -255 -17 -252
rect 16 -255 28 -252
rect 76 -252 79 -249
rect -97 -260 -85 -258
rect -92 -261 -85 -260
rect -88 -264 -85 -261
rect -80 -264 -77 -257
rect -69 -262 -63 -259
rect -22 -263 -19 -255
rect -52 -266 -19 -263
rect 18 -263 21 -255
rect 62 -262 68 -259
rect 18 -266 51 -263
rect 76 -264 79 -257
rect -52 -269 -49 -266
rect -65 -271 -49 -269
rect -68 -272 -49 -271
rect 48 -269 51 -266
rect 84 -258 87 -251
rect 84 -260 96 -258
rect 84 -261 91 -260
rect 84 -264 87 -261
rect 125 -264 128 -257
rect 191 -250 194 -240
rect 209 -244 216 -240
rect 224 -249 227 -205
rect 302 -206 365 -203
rect 271 -217 274 -215
rect 257 -229 258 -224
rect 263 -227 264 -224
rect 263 -229 290 -227
rect 257 -230 290 -229
rect 257 -231 264 -230
rect 268 -237 271 -230
rect 206 -252 219 -249
rect 226 -253 227 -249
rect 231 -240 280 -237
rect 231 -250 234 -240
rect 133 -258 136 -255
rect 184 -261 196 -258
rect 229 -261 241 -258
rect 289 -258 292 -255
rect 116 -266 128 -264
rect 48 -271 64 -269
rect 48 -272 67 -271
rect -68 -274 -62 -272
rect -65 -277 -62 -274
rect -79 -280 -62 -277
rect 61 -274 67 -272
rect 121 -267 128 -266
rect 125 -270 128 -267
rect 133 -270 136 -263
rect 144 -268 150 -265
rect 191 -269 194 -261
rect 161 -272 194 -269
rect 231 -269 234 -261
rect 275 -268 281 -265
rect 231 -272 264 -269
rect 289 -270 292 -263
rect 61 -277 64 -274
rect 161 -275 164 -272
rect 61 -280 78 -277
rect 148 -277 164 -275
rect 145 -278 164 -277
rect 261 -275 264 -272
rect 297 -264 300 -257
rect 297 -266 309 -264
rect 297 -267 304 -266
rect 297 -270 300 -267
rect 261 -277 277 -275
rect 261 -278 280 -277
rect 145 -280 151 -278
rect 148 -283 151 -280
rect 134 -286 151 -283
rect 274 -280 280 -278
rect 274 -283 277 -280
rect 274 -286 291 -283
<< m2contact >>
rect 365 -76 370 -71
rect 346 -85 351 -80
rect 282 -120 287 -115
rect 291 -122 296 -117
rect -46 -170 -40 -165
rect -55 -181 -50 -176
rect -5 -171 0 -166
rect 28 -177 33 -172
rect -39 -189 -34 -184
rect -5 -187 0 -182
rect -63 -216 -58 -211
rect -9 -239 -4 -234
rect 3 -239 8 -234
rect 22 -200 27 -195
rect 60 -182 65 -177
rect 168 -176 173 -171
rect 110 -185 115 -180
rect 52 -199 57 -194
rect 94 -200 99 -195
rect 157 -203 162 -198
rect 174 -186 179 -181
rect 208 -177 213 -172
rect 249 -175 254 -170
rect 353 -181 358 -176
rect 174 -195 179 -190
rect 208 -193 213 -188
rect 244 -190 249 -185
rect 57 -216 62 -211
rect 115 -213 120 -208
rect 354 -192 359 -187
rect 150 -222 155 -217
rect -81 -257 -76 -252
rect 75 -257 80 -252
rect 204 -245 209 -240
rect 216 -245 221 -240
rect 270 -222 275 -217
rect 132 -263 137 -258
rect 288 -263 293 -258
<< pdm12contact >>
rect -49 -247 -44 -242
rect 43 -247 48 -242
rect 164 -253 169 -248
rect 256 -253 261 -248
<< metal2 >>
rect 348 -75 365 -72
rect 348 -80 351 -75
rect 200 -111 223 -108
rect 200 -132 203 -111
rect 220 -117 223 -111
rect 220 -120 282 -117
rect 296 -121 358 -118
rect 111 -135 203 -132
rect 111 -157 114 -135
rect 250 -136 309 -133
rect -54 -160 114 -157
rect -54 -176 -51 -160
rect -40 -169 -5 -166
rect -46 -201 -43 -170
rect 29 -178 33 -177
rect 29 -181 60 -178
rect -34 -187 -5 -184
rect 111 -180 114 -160
rect 160 -182 163 -149
rect 250 -170 253 -136
rect 173 -175 208 -172
rect 355 -176 358 -121
rect 318 -180 353 -177
rect 160 -185 174 -182
rect 27 -199 52 -196
rect 179 -193 208 -190
rect 318 -186 321 -180
rect 249 -189 321 -186
rect 359 -191 377 -187
rect 99 -199 115 -196
rect -54 -204 -43 -201
rect -54 -212 -51 -204
rect -58 -215 -51 -212
rect -101 -253 -98 -225
rect -101 -256 -81 -253
rect -62 -258 -59 -216
rect 112 -212 115 -199
rect 162 -202 180 -199
rect 177 -210 180 -202
rect 177 -213 274 -210
rect -48 -230 -13 -227
rect -48 -242 -45 -230
rect -16 -235 -13 -230
rect 12 -230 47 -227
rect -16 -238 -9 -235
rect 12 -235 15 -230
rect 8 -238 15 -235
rect 44 -242 47 -230
rect 58 -258 61 -216
rect 271 -217 274 -213
rect 80 -256 103 -253
rect 100 -282 103 -256
rect 112 -259 115 -231
rect 112 -262 132 -259
rect 151 -264 154 -222
rect 165 -236 200 -233
rect 165 -248 168 -236
rect 197 -241 200 -236
rect 225 -236 260 -233
rect 197 -244 204 -241
rect 225 -241 228 -236
rect 221 -244 228 -241
rect 257 -248 260 -236
rect 271 -264 274 -222
rect 293 -262 316 -259
rect 313 -288 316 -262
<< m3contact >>
rect 159 -149 164 -144
rect 29 -186 34 -181
rect 309 -137 314 -132
rect 377 -192 382 -187
rect -102 -225 -97 -220
rect 111 -231 116 -226
<< m123contact >>
rect -3 -115 2 -110
rect 210 -121 215 -116
rect 264 -112 269 -107
rect 364 -121 369 -116
rect 308 -175 313 -170
rect 406 -141 411 -136
rect -3 -218 2 -213
rect 265 -204 270 -199
rect 45 -223 50 -218
rect -97 -265 -92 -260
rect -63 -263 -58 -258
rect 57 -263 62 -258
rect 91 -265 96 -260
rect 210 -224 215 -219
rect 258 -229 263 -224
rect 116 -271 121 -266
rect 150 -269 155 -264
rect 270 -269 275 -264
rect 304 -271 309 -266
<< metal3 >>
rect 255 -103 364 -100
rect 195 -107 228 -104
rect -2 -213 1 -115
rect 195 -127 198 -107
rect 225 -112 228 -107
rect 255 -112 258 -103
rect 225 -115 258 -112
rect 160 -130 198 -127
rect 160 -143 163 -130
rect 158 -144 165 -143
rect 158 -149 159 -144
rect 164 -149 165 -144
rect 158 -150 165 -149
rect 28 -181 35 -180
rect 28 -186 29 -181
rect 34 -186 35 -181
rect 28 -187 35 -186
rect 29 -203 33 -187
rect 153 -203 157 -169
rect 29 -207 157 -203
rect -103 -220 -96 -219
rect -103 -225 -102 -220
rect -97 -222 -96 -220
rect 44 -222 45 -218
rect -97 -223 45 -222
rect 50 -223 51 -218
rect 211 -219 214 -121
rect 265 -199 268 -112
rect 361 -120 364 -103
rect 308 -132 315 -131
rect 308 -137 309 -132
rect 314 -133 315 -132
rect 314 -136 407 -133
rect 314 -137 315 -136
rect 308 -138 315 -137
rect 404 -139 406 -136
rect -97 -225 51 -223
rect -103 -226 -96 -225
rect 110 -226 117 -225
rect 110 -231 111 -226
rect 116 -228 117 -226
rect 257 -228 258 -224
rect 116 -229 258 -228
rect 263 -229 264 -224
rect 116 -231 264 -229
rect 110 -232 117 -231
rect 309 -245 312 -175
rect 377 -186 381 -169
rect 376 -187 383 -186
rect 376 -192 377 -187
rect 382 -192 383 -187
rect 376 -193 383 -192
rect 174 -248 312 -245
rect -95 -260 -63 -259
rect -92 -262 -63 -260
rect 62 -260 94 -259
rect 62 -262 91 -260
rect 92 -278 95 -265
rect 118 -266 150 -265
rect 121 -268 150 -266
rect 174 -278 177 -248
rect 275 -266 307 -265
rect 275 -268 304 -266
rect 92 -281 177 -278
<< m4contact >>
rect 153 -169 158 -164
rect 377 -169 382 -164
<< metal4 >>
rect 158 -169 377 -165
<< labels >>
rlabel metal1 -1 -236 -1 -236 3 vdd
rlabel metal1 -1 -244 -1 -244 3 gnd
rlabel metal1 -15 -136 -15 -136 5 vdd
rlabel metal1 14 -197 14 -197 1 gnd
rlabel metal1 4 -116 4 -115 5 vdd
rlabel metal1 138 -182 144 -179 7 c1
rlabel metal1 131 -211 131 -211 1 gnd
rlabel metal1 122 -138 122 -138 5 vdd
rlabel m2contact 61 -179 65 -178 1 p0_inv
rlabel metal1 105 -175 107 -172 1 temp100
rlabel metal1 68 -116 68 -115 5 vdd
rlabel metal1 78 -197 78 -197 1 gnd
rlabel metal1 53 -153 55 -150 1 c0_inv
rlabel metal1 38 -154 40 -152 3 c0
rlabel metal1 44 -173 44 -173 1 gnd
rlabel metal1 43 -115 43 -115 5 vdd
rlabel m2contact 59 -214 60 -214 1 c0
rlabel metal2 101 -282 102 -280 1 s0
rlabel metal2 -100 -255 -96 -253 3 mid_s0
rlabel metal1 -8 -174 3 -171 1 a0
rlabel metal1 -8 -181 3 -178 1 b0
rlabel metal1 -37 -180 -31 -177 1 g0_inv
rlabel metal1 25 -176 30 -173 1 p0_inv
rlabel m2contact 111 -183 115 -181 1 g0_inv
rlabel metal1 212 -242 212 -242 3 vdd
rlabel metal1 212 -250 212 -250 3 gnd
rlabel metal1 198 -142 198 -142 5 vdd
rlabel metal1 227 -203 227 -203 1 gnd
rlabel metal1 217 -122 217 -121 5 vdd
rlabel metal2 113 -260 113 -260 1 mid_s1
rlabel metal2 314 -288 315 -286 8 s1
rlabel metal1 176 -186 182 -183 1 g1_inv
rlabel metal1 238 -182 243 -179 1 p1_inv
rlabel metal1 205 -180 216 -177 1 a1
rlabel metal1 205 -187 216 -184 1 b1
rlabel metal1 272 -218 274 -215 1 c1
rlabel metal1 350 -123 350 -122 5 vdd
rlabel metal1 340 -204 340 -204 1 gnd
rlabel metal1 351 -181 355 -179 7 p1_inv
rlabel metal1 352 -187 357 -185 7 p0_inv
rlabel metal1 324 -183 328 -181 3 temp101
rlabel metal1 294 -129 294 -129 5 vdd
rlabel metal1 285 -202 285 -202 1 gnd
rlabel metal1 301 -173 305 -172 1 c0
rlabel metal1 257 -172 259 -170 1 temp102
rlabel metal1 268 -100 268 -100 3 gnd
rlabel metal1 349 -110 350 -110 7 vdd
rlabel space 285 -116 288 -113 1 g0_inv
rlabel metal1 290 -74 293 -71 1 temp103
rlabel metal1 377 -75 377 -75 5 vdd
rlabel metal1 386 -148 386 -148 1 gnd
rlabel metal1 393 -119 399 -116 7 temp104
rlabel metal1 415 -75 415 -74 5 vdd
rlabel metal1 425 -156 425 -156 1 gnd
rlabel metal1 452 -134 454 -132 1 c2
rlabel m123contact 365 -119 365 -119 1 g1_inv
<< end >>
