magic
tech scmos
timestamp 1731612933
<< nwell >>
rect -203 344 -126 366
rect -86 360 -54 379
rect -221 334 -126 344
rect -108 354 -54 360
rect -221 314 -169 334
rect -108 326 -56 354
rect -221 312 -197 314
rect -389 279 -357 298
rect -389 273 -335 279
rect -387 245 -335 273
rect -317 263 -240 285
rect -118 266 -84 318
rect -67 306 -33 312
rect -67 280 -11 306
rect -36 274 -11 280
rect -317 253 -222 263
rect -410 225 -376 231
rect -432 199 -376 225
rect -432 193 -407 199
rect -359 185 -325 237
rect -274 233 -222 253
rect -246 231 -222 233
rect -552 144 -494 166
rect -292 157 -231 189
rect -552 134 -445 144
rect -623 93 -562 125
rect -528 114 -445 134
rect -500 112 -445 114
rect -429 105 -368 137
rect -268 40 -207 41
rect -577 37 -516 38
rect -417 37 -356 38
rect -577 26 -479 37
rect -417 26 -319 37
rect -268 29 -170 40
rect -577 6 -445 26
rect -417 6 -285 26
rect -268 9 -136 29
rect -513 -6 -445 6
rect -353 -6 -285 6
rect -204 -3 -136 9
rect -513 -15 -479 -6
rect -353 -15 -319 -6
rect -204 -12 -170 -3
<< ntransistor >>
rect -48 365 -38 367
rect -44 347 -34 349
rect -44 337 -34 339
rect -210 296 -208 306
rect -149 302 -147 322
rect -139 302 -137 322
rect -192 292 -190 302
rect -182 292 -180 302
rect -405 284 -395 286
rect -409 266 -399 268
rect -409 256 -399 258
rect -306 221 -304 241
rect -296 221 -294 241
rect -107 244 -105 254
rect -97 244 -95 254
rect -56 248 -54 268
rect -46 248 -44 268
rect -25 258 -23 268
rect -263 211 -261 221
rect -253 211 -251 221
rect -235 215 -233 225
rect -420 177 -418 187
rect -399 167 -397 187
rect -389 167 -387 187
rect -348 163 -346 173
rect -338 163 -336 173
rect -541 118 -539 128
rect -281 140 -279 150
rect -272 140 -270 150
rect -244 141 -242 151
rect -517 92 -515 102
rect -507 92 -505 102
rect -489 96 -487 106
rect -612 76 -610 86
rect -603 76 -601 86
rect -575 77 -573 87
rect -468 80 -466 100
rect -458 80 -456 100
rect -418 88 -416 98
rect -409 88 -407 98
rect -381 89 -379 99
rect -566 45 -564 55
rect -557 45 -555 55
rect -529 44 -527 54
rect -502 49 -500 59
rect -492 49 -490 59
rect -468 38 -466 58
rect -458 38 -456 58
rect -406 45 -404 55
rect -397 45 -395 55
rect -369 44 -367 54
rect -342 49 -340 59
rect -332 49 -330 59
rect -308 38 -306 58
rect -298 38 -296 58
rect -257 48 -255 58
rect -248 48 -246 58
rect -220 47 -218 57
rect -193 52 -191 62
rect -183 52 -181 62
rect -159 41 -157 61
rect -149 41 -147 61
<< ptransistor >>
rect -80 365 -60 367
rect -210 318 -208 338
rect -192 320 -190 360
rect -182 320 -180 360
rect -149 340 -147 360
rect -139 340 -137 360
rect -102 347 -62 349
rect -102 337 -62 339
rect -383 284 -363 286
rect -381 266 -341 268
rect -306 259 -304 279
rect -296 259 -294 279
rect -381 256 -341 258
rect -420 199 -418 219
rect -399 205 -397 225
rect -389 205 -387 225
rect -348 191 -346 231
rect -338 191 -336 231
rect -263 239 -261 279
rect -253 239 -251 279
rect -107 272 -105 312
rect -97 272 -95 312
rect -56 286 -54 306
rect -46 286 -44 306
rect -235 237 -233 257
rect -25 280 -23 300
rect -281 163 -279 183
rect -272 163 -270 183
rect -244 163 -242 183
rect -541 140 -539 160
rect -612 99 -610 119
rect -603 99 -601 119
rect -575 99 -573 119
rect -517 120 -515 160
rect -507 120 -505 160
rect -489 118 -487 138
rect -468 118 -466 138
rect -458 118 -456 138
rect -418 111 -416 131
rect -409 111 -407 131
rect -381 111 -379 131
rect -566 12 -564 32
rect -557 12 -555 32
rect -529 12 -527 32
rect -502 -9 -500 31
rect -492 -9 -490 31
rect -468 0 -466 20
rect -458 0 -456 20
rect -406 12 -404 32
rect -397 12 -395 32
rect -369 12 -367 32
rect -342 -9 -340 31
rect -332 -9 -330 31
rect -308 0 -306 20
rect -298 0 -296 20
rect -257 15 -255 35
rect -248 15 -246 35
rect -220 15 -218 35
rect -193 -6 -191 34
rect -183 -6 -181 34
rect -159 3 -157 23
rect -149 3 -147 23
<< ndiffusion >>
rect -44 368 -38 372
rect -48 367 -38 368
rect -48 364 -38 365
rect -48 360 -42 364
rect -44 350 -38 354
rect -44 349 -34 350
rect -44 345 -34 347
rect -40 341 -34 345
rect -44 339 -34 341
rect -44 336 -34 337
rect -44 332 -38 336
rect -211 302 -210 306
rect -215 296 -210 302
rect -208 300 -203 306
rect -150 318 -149 322
rect -154 302 -149 318
rect -147 302 -139 322
rect -137 306 -132 322
rect -137 302 -136 306
rect -208 296 -207 300
rect -197 296 -192 302
rect -193 292 -192 296
rect -190 298 -188 302
rect -184 298 -182 302
rect -190 292 -182 298
rect -180 296 -175 302
rect -180 292 -179 296
rect -405 287 -399 291
rect -405 286 -395 287
rect -405 283 -395 284
rect -401 279 -395 283
rect -405 269 -399 273
rect -409 268 -399 269
rect -409 264 -399 266
rect -409 260 -403 264
rect -409 258 -399 260
rect -409 255 -399 256
rect -405 251 -399 255
rect -311 225 -306 241
rect -307 221 -306 225
rect -304 221 -296 241
rect -294 237 -293 241
rect -294 221 -289 237
rect -112 248 -107 254
rect -108 244 -107 248
rect -105 250 -103 254
rect -99 250 -97 254
rect -105 244 -97 250
rect -95 248 -90 254
rect -61 252 -56 268
rect -57 248 -56 252
rect -54 248 -46 268
rect -44 264 -43 268
rect -44 248 -39 264
rect -30 262 -25 268
rect -26 258 -25 262
rect -23 264 -22 268
rect -23 258 -18 264
rect -95 244 -94 248
rect -268 215 -263 221
rect -264 211 -263 215
rect -261 217 -259 221
rect -255 217 -253 221
rect -261 211 -253 217
rect -251 215 -246 221
rect -240 219 -235 225
rect -236 215 -235 219
rect -233 221 -232 225
rect -233 215 -228 221
rect -251 211 -250 215
rect -421 183 -420 187
rect -425 177 -420 183
rect -418 181 -413 187
rect -418 177 -417 181
rect -400 183 -399 187
rect -404 167 -399 183
rect -397 167 -389 187
rect -387 171 -382 187
rect -387 167 -386 171
rect -353 167 -348 173
rect -349 163 -348 167
rect -346 169 -344 173
rect -340 169 -338 173
rect -346 163 -338 169
rect -336 167 -331 173
rect -336 163 -335 167
rect -546 122 -541 128
rect -542 118 -541 122
rect -539 124 -538 128
rect -539 118 -534 124
rect -282 146 -281 150
rect -286 140 -281 146
rect -279 146 -277 150
rect -273 146 -272 150
rect -279 140 -272 146
rect -270 144 -265 150
rect -270 140 -269 144
rect -249 145 -244 151
rect -245 141 -244 145
rect -242 145 -237 151
rect -242 141 -241 145
rect -522 96 -517 102
rect -518 92 -517 96
rect -515 98 -513 102
rect -509 98 -507 102
rect -515 92 -507 98
rect -505 96 -500 102
rect -494 100 -489 106
rect -490 96 -489 100
rect -487 102 -486 106
rect -487 96 -482 102
rect -505 92 -504 96
rect -613 82 -612 86
rect -617 76 -612 82
rect -610 82 -608 86
rect -604 82 -603 86
rect -610 76 -603 82
rect -601 80 -596 86
rect -601 76 -600 80
rect -580 81 -575 87
rect -576 77 -575 81
rect -573 81 -568 87
rect -573 77 -572 81
rect -473 84 -468 100
rect -469 80 -468 84
rect -466 80 -458 100
rect -456 96 -455 100
rect -456 80 -451 96
rect -419 94 -418 98
rect -423 88 -418 94
rect -416 94 -414 98
rect -410 94 -409 98
rect -416 88 -409 94
rect -407 92 -402 98
rect -407 88 -406 92
rect -386 93 -381 99
rect -382 89 -381 93
rect -379 93 -374 99
rect -379 89 -378 93
rect -571 49 -566 55
rect -567 45 -566 49
rect -564 49 -557 55
rect -564 45 -562 49
rect -558 45 -557 49
rect -555 51 -554 55
rect -503 55 -502 59
rect -555 45 -550 51
rect -530 50 -529 54
rect -534 44 -529 50
rect -527 50 -526 54
rect -527 44 -522 50
rect -507 49 -502 55
rect -500 53 -492 59
rect -500 49 -498 53
rect -494 49 -492 53
rect -490 55 -489 59
rect -490 49 -485 55
rect -469 54 -468 58
rect -473 38 -468 54
rect -466 38 -458 58
rect -456 42 -451 58
rect -411 49 -406 55
rect -407 45 -406 49
rect -404 49 -397 55
rect -404 45 -402 49
rect -398 45 -397 49
rect -395 51 -394 55
rect -343 55 -342 59
rect -395 45 -390 51
rect -370 50 -369 54
rect -456 38 -455 42
rect -374 44 -369 50
rect -367 50 -366 54
rect -367 44 -362 50
rect -347 49 -342 55
rect -340 53 -332 59
rect -340 49 -338 53
rect -334 49 -332 53
rect -330 55 -329 59
rect -330 49 -325 55
rect -309 54 -308 58
rect -313 38 -308 54
rect -306 38 -298 58
rect -296 42 -291 58
rect -262 52 -257 58
rect -258 48 -257 52
rect -255 52 -248 58
rect -255 48 -253 52
rect -249 48 -248 52
rect -246 54 -245 58
rect -194 58 -193 62
rect -246 48 -241 54
rect -221 53 -220 57
rect -296 38 -295 42
rect -225 47 -220 53
rect -218 53 -217 57
rect -218 47 -213 53
rect -198 52 -193 58
rect -191 56 -183 62
rect -191 52 -189 56
rect -185 52 -183 56
rect -181 58 -180 62
rect -181 52 -176 58
rect -160 57 -159 61
rect -164 41 -159 57
rect -157 41 -149 61
rect -147 45 -142 61
rect -147 41 -146 45
<< pdiffusion >>
rect -80 368 -64 372
rect -80 367 -60 368
rect -80 364 -60 365
rect -76 360 -60 364
rect -215 322 -210 338
rect -211 318 -210 322
rect -208 334 -207 338
rect -208 318 -203 334
rect -197 324 -192 360
rect -193 320 -192 324
rect -190 320 -182 360
rect -180 356 -179 360
rect -180 320 -175 356
rect -150 356 -149 360
rect -154 340 -149 356
rect -147 344 -139 360
rect -147 340 -145 344
rect -141 340 -139 344
rect -137 356 -136 360
rect -137 340 -132 356
rect -102 350 -66 354
rect -102 349 -62 350
rect -102 339 -62 347
rect -102 336 -62 337
rect -98 332 -62 336
rect -108 308 -107 312
rect -379 287 -363 291
rect -383 286 -363 287
rect -383 283 -363 284
rect -383 279 -367 283
rect -307 275 -306 279
rect -377 269 -341 273
rect -381 268 -341 269
rect -381 258 -341 266
rect -311 259 -306 275
rect -304 263 -296 279
rect -304 259 -302 263
rect -298 259 -296 263
rect -294 275 -293 279
rect -294 259 -289 275
rect -264 275 -263 279
rect -381 255 -341 256
rect -381 251 -345 255
rect -400 221 -399 225
rect -425 203 -420 219
rect -421 199 -420 203
rect -418 215 -417 219
rect -418 199 -413 215
rect -404 205 -399 221
rect -397 209 -389 225
rect -397 205 -395 209
rect -391 205 -389 209
rect -387 221 -386 225
rect -387 205 -382 221
rect -353 195 -348 231
rect -349 191 -348 195
rect -346 191 -338 231
rect -336 227 -335 231
rect -336 191 -331 227
rect -268 239 -263 275
rect -261 239 -253 279
rect -251 243 -246 279
rect -112 272 -107 308
rect -105 272 -97 312
rect -95 276 -90 312
rect -57 302 -56 306
rect -61 286 -56 302
rect -54 290 -46 306
rect -54 286 -52 290
rect -48 286 -46 290
rect -44 302 -43 306
rect -44 286 -39 302
rect -26 296 -25 300
rect -95 272 -94 276
rect -251 239 -250 243
rect -236 253 -235 257
rect -240 237 -235 253
rect -233 241 -228 257
rect -30 280 -25 296
rect -23 284 -18 300
rect -23 280 -22 284
rect -233 237 -232 241
rect -286 167 -281 183
rect -282 163 -281 167
rect -279 169 -272 183
rect -279 165 -277 169
rect -273 165 -272 169
rect -279 163 -272 165
rect -270 179 -269 183
rect -270 163 -265 179
rect -245 179 -244 183
rect -249 163 -244 179
rect -242 167 -237 183
rect -242 163 -241 167
rect -542 156 -541 160
rect -546 140 -541 156
rect -539 144 -534 160
rect -539 140 -538 144
rect -518 156 -517 160
rect -617 103 -612 119
rect -613 99 -612 103
rect -610 105 -603 119
rect -610 101 -608 105
rect -604 101 -603 105
rect -610 99 -603 101
rect -601 115 -600 119
rect -601 99 -596 115
rect -576 115 -575 119
rect -580 99 -575 115
rect -573 103 -568 119
rect -522 120 -517 156
rect -515 120 -507 160
rect -505 124 -500 160
rect -505 120 -504 124
rect -490 134 -489 138
rect -573 99 -572 103
rect -494 118 -489 134
rect -487 122 -482 138
rect -487 118 -486 122
rect -469 134 -468 138
rect -473 118 -468 134
rect -466 122 -458 138
rect -466 118 -464 122
rect -460 118 -458 122
rect -456 134 -455 138
rect -456 118 -451 134
rect -423 115 -418 131
rect -419 111 -418 115
rect -416 117 -409 131
rect -416 113 -414 117
rect -410 113 -409 117
rect -416 111 -409 113
rect -407 127 -406 131
rect -407 111 -402 127
rect -382 127 -381 131
rect -386 111 -381 127
rect -379 115 -374 131
rect -379 111 -378 115
rect -567 28 -566 32
rect -571 12 -566 28
rect -564 30 -557 32
rect -564 26 -562 30
rect -558 26 -557 30
rect -564 12 -557 26
rect -555 16 -550 32
rect -555 12 -554 16
rect -534 16 -529 32
rect -530 12 -529 16
rect -527 28 -526 32
rect -527 12 -522 28
rect -507 -5 -502 31
rect -503 -9 -502 -5
rect -500 -9 -492 31
rect -490 27 -489 31
rect -490 -9 -485 27
rect -407 28 -406 32
rect -473 4 -468 20
rect -469 0 -468 4
rect -466 16 -464 20
rect -460 16 -458 20
rect -466 0 -458 16
rect -456 4 -451 20
rect -411 12 -406 28
rect -404 30 -397 32
rect -404 26 -402 30
rect -398 26 -397 30
rect -404 12 -397 26
rect -395 16 -390 32
rect -395 12 -394 16
rect -374 16 -369 32
rect -370 12 -369 16
rect -367 28 -366 32
rect -367 12 -362 28
rect -456 0 -455 4
rect -347 -5 -342 31
rect -343 -9 -342 -5
rect -340 -9 -332 31
rect -330 27 -329 31
rect -330 -9 -325 27
rect -258 31 -257 35
rect -313 4 -308 20
rect -309 0 -308 4
rect -306 16 -304 20
rect -300 16 -298 20
rect -306 0 -298 16
rect -296 4 -291 20
rect -262 15 -257 31
rect -255 33 -248 35
rect -255 29 -253 33
rect -249 29 -248 33
rect -255 15 -248 29
rect -246 19 -241 35
rect -246 15 -245 19
rect -225 19 -220 35
rect -221 15 -220 19
rect -218 31 -217 35
rect -218 15 -213 31
rect -296 0 -295 4
rect -198 -2 -193 34
rect -194 -6 -193 -2
rect -191 -6 -183 34
rect -181 30 -180 34
rect -181 -6 -176 30
rect -164 7 -159 23
rect -160 3 -159 7
rect -157 19 -155 23
rect -151 19 -149 23
rect -157 3 -149 19
rect -147 7 -142 23
rect -147 3 -146 7
<< ndcontact >>
rect -48 368 -44 372
rect -42 360 -38 364
rect -38 350 -34 354
rect -44 341 -40 345
rect -38 332 -34 336
rect -215 302 -211 306
rect -154 318 -150 322
rect -136 302 -132 306
rect -207 296 -203 300
rect -197 292 -193 296
rect -188 298 -184 302
rect -179 292 -175 296
rect -399 287 -395 291
rect -405 279 -401 283
rect -409 269 -405 273
rect -403 260 -399 264
rect -409 251 -405 255
rect -311 221 -307 225
rect -293 237 -289 241
rect -112 244 -108 248
rect -103 250 -99 254
rect -61 248 -57 252
rect -43 264 -39 268
rect -30 258 -26 262
rect -22 264 -18 268
rect -94 244 -90 248
rect -268 211 -264 215
rect -259 217 -255 221
rect -240 215 -236 219
rect -232 221 -228 225
rect -250 211 -246 215
rect -425 183 -421 187
rect -417 177 -413 181
rect -404 183 -400 187
rect -386 167 -382 171
rect -353 163 -349 167
rect -344 169 -340 173
rect -335 163 -331 167
rect -546 118 -542 122
rect -538 124 -534 128
rect -286 146 -282 150
rect -277 146 -273 150
rect -269 140 -265 144
rect -249 141 -245 145
rect -241 141 -237 145
rect -522 92 -518 96
rect -513 98 -509 102
rect -494 96 -490 100
rect -486 102 -482 106
rect -504 92 -500 96
rect -617 82 -613 86
rect -608 82 -604 86
rect -600 76 -596 80
rect -580 77 -576 81
rect -572 77 -568 81
rect -473 80 -469 84
rect -455 96 -451 100
rect -423 94 -419 98
rect -414 94 -410 98
rect -406 88 -402 92
rect -386 89 -382 93
rect -378 89 -374 93
rect -571 45 -567 49
rect -562 45 -558 49
rect -554 51 -550 55
rect -507 55 -503 59
rect -534 50 -530 54
rect -526 50 -522 54
rect -498 49 -494 53
rect -489 55 -485 59
rect -473 54 -469 58
rect -411 45 -407 49
rect -402 45 -398 49
rect -394 51 -390 55
rect -347 55 -343 59
rect -374 50 -370 54
rect -455 38 -451 42
rect -366 50 -362 54
rect -338 49 -334 53
rect -329 55 -325 59
rect -313 54 -309 58
rect -262 48 -258 52
rect -253 48 -249 52
rect -245 54 -241 58
rect -198 58 -194 62
rect -225 53 -221 57
rect -295 38 -291 42
rect -217 53 -213 57
rect -189 52 -185 56
rect -180 58 -176 62
rect -164 57 -160 61
rect -146 41 -142 45
<< pdcontact >>
rect -64 368 -60 372
rect -80 360 -76 364
rect -215 318 -211 322
rect -207 334 -203 338
rect -197 320 -193 324
rect -179 356 -175 360
rect -154 356 -150 360
rect -145 340 -141 344
rect -136 356 -132 360
rect -66 350 -62 354
rect -102 332 -98 336
rect -112 308 -108 312
rect -383 287 -379 291
rect -367 279 -363 283
rect -311 275 -307 279
rect -381 269 -377 273
rect -302 259 -298 263
rect -293 275 -289 279
rect -268 275 -264 279
rect -345 251 -341 255
rect -404 221 -400 225
rect -425 199 -421 203
rect -417 215 -413 219
rect -395 205 -391 209
rect -386 221 -382 225
rect -353 191 -349 195
rect -335 227 -331 231
rect -61 302 -57 306
rect -52 286 -48 290
rect -43 302 -39 306
rect -30 296 -26 300
rect -94 272 -90 276
rect -250 239 -246 243
rect -240 253 -236 257
rect -22 280 -18 284
rect -232 237 -228 241
rect -286 163 -282 167
rect -277 165 -273 169
rect -269 179 -265 183
rect -249 179 -245 183
rect -241 163 -237 167
rect -546 156 -542 160
rect -538 140 -534 144
rect -522 156 -518 160
rect -617 99 -613 103
rect -608 101 -604 105
rect -600 115 -596 119
rect -580 115 -576 119
rect -504 120 -500 124
rect -494 134 -490 138
rect -572 99 -568 103
rect -486 118 -482 122
rect -473 134 -469 138
rect -464 118 -460 122
rect -455 134 -451 138
rect -423 111 -419 115
rect -414 113 -410 117
rect -406 127 -402 131
rect -386 127 -382 131
rect -378 111 -374 115
rect -571 28 -567 32
rect -562 26 -558 30
rect -554 12 -550 16
rect -534 12 -530 16
rect -526 28 -522 32
rect -507 -9 -503 -5
rect -489 27 -485 31
rect -411 28 -407 32
rect -473 0 -469 4
rect -464 16 -460 20
rect -402 26 -398 30
rect -394 12 -390 16
rect -374 12 -370 16
rect -366 28 -362 32
rect -455 0 -451 4
rect -347 -9 -343 -5
rect -329 27 -325 31
rect -262 31 -258 35
rect -313 0 -309 4
rect -304 16 -300 20
rect -253 29 -249 33
rect -245 15 -241 19
rect -225 15 -221 19
rect -217 31 -213 35
rect -295 0 -291 4
rect -198 -6 -194 -2
rect -180 30 -176 34
rect -164 3 -160 7
rect -155 19 -151 23
rect -146 3 -142 7
<< polysilicon >>
rect -83 365 -80 367
rect -60 365 -48 367
rect -38 365 -35 367
rect -192 360 -190 363
rect -182 360 -180 363
rect -149 360 -147 364
rect -139 360 -137 364
rect -210 338 -208 341
rect -105 347 -102 349
rect -62 347 -44 349
rect -34 347 -31 349
rect -149 322 -147 340
rect -139 322 -137 340
rect -105 337 -102 339
rect -62 337 -44 339
rect -34 337 -31 339
rect -210 306 -208 318
rect -192 302 -190 320
rect -182 302 -180 320
rect -107 312 -105 315
rect -97 312 -95 315
rect -210 293 -208 296
rect -149 298 -147 302
rect -139 298 -137 302
rect -192 289 -190 292
rect -182 289 -180 292
rect -408 284 -405 286
rect -395 284 -383 286
rect -363 284 -360 286
rect -306 279 -304 283
rect -296 279 -294 283
rect -263 279 -261 282
rect -253 279 -251 282
rect -412 266 -409 268
rect -399 266 -381 268
rect -341 266 -338 268
rect -412 256 -409 258
rect -399 256 -381 258
rect -341 256 -338 258
rect -306 241 -304 259
rect -296 241 -294 259
rect -348 231 -346 234
rect -338 231 -336 234
rect -399 225 -397 229
rect -389 225 -387 229
rect -420 219 -418 223
rect -420 187 -418 199
rect -399 187 -397 205
rect -389 187 -387 205
rect -56 306 -54 310
rect -46 306 -44 310
rect -25 300 -23 304
rect -235 257 -233 260
rect -263 221 -261 239
rect -253 221 -251 239
rect -107 254 -105 272
rect -97 254 -95 272
rect -56 268 -54 286
rect -46 268 -44 286
rect -25 268 -23 280
rect -25 254 -23 258
rect -56 244 -54 248
rect -46 244 -44 248
rect -107 241 -105 244
rect -97 241 -95 244
rect -235 225 -233 237
rect -306 217 -304 221
rect -296 217 -294 221
rect -235 212 -233 215
rect -263 208 -261 211
rect -253 208 -251 211
rect -420 173 -418 177
rect -348 173 -346 191
rect -338 173 -336 191
rect -281 183 -279 195
rect -272 183 -270 186
rect -244 183 -242 187
rect -541 160 -539 164
rect -399 163 -397 167
rect -389 163 -387 167
rect -517 160 -515 163
rect -507 160 -505 163
rect -348 160 -346 163
rect -338 160 -336 163
rect -612 119 -610 131
rect -541 128 -539 140
rect -603 119 -601 122
rect -575 119 -573 123
rect -281 157 -279 163
rect -281 150 -279 154
rect -272 150 -270 163
rect -244 151 -242 163
rect -489 138 -487 141
rect -468 138 -466 142
rect -458 138 -456 142
rect -541 114 -539 118
rect -517 102 -515 120
rect -507 102 -505 120
rect -418 131 -416 143
rect -281 138 -279 140
rect -409 131 -407 134
rect -381 131 -379 135
rect -281 134 -280 138
rect -272 137 -270 140
rect -244 137 -242 141
rect -281 133 -279 134
rect -489 106 -487 118
rect -612 93 -610 99
rect -612 86 -610 90
rect -603 86 -601 99
rect -575 87 -573 99
rect -468 100 -466 118
rect -458 100 -456 118
rect -418 105 -416 111
rect -489 93 -487 96
rect -517 89 -515 92
rect -507 89 -505 92
rect -418 98 -416 102
rect -409 98 -407 111
rect -381 99 -379 111
rect -418 86 -416 88
rect -418 82 -417 86
rect -409 85 -407 88
rect -381 85 -379 89
rect -418 81 -416 82
rect -612 74 -610 76
rect -612 70 -611 74
rect -603 73 -601 76
rect -575 73 -573 77
rect -468 76 -466 80
rect -458 76 -456 80
rect -612 69 -610 70
rect -257 64 -255 65
rect -566 61 -564 62
rect -566 57 -565 61
rect -502 59 -500 62
rect -492 59 -490 62
rect -566 55 -564 57
rect -557 55 -555 58
rect -529 54 -527 58
rect -566 41 -564 45
rect -566 32 -564 38
rect -557 32 -555 45
rect -468 58 -466 62
rect -458 58 -456 62
rect -406 61 -404 62
rect -529 32 -527 44
rect -502 31 -500 49
rect -492 31 -490 49
rect -406 57 -405 61
rect -342 59 -340 62
rect -332 59 -330 62
rect -406 55 -404 57
rect -397 55 -395 58
rect -369 54 -367 58
rect -406 41 -404 45
rect -566 0 -564 12
rect -557 9 -555 12
rect -529 8 -527 12
rect -468 20 -466 38
rect -458 20 -456 38
rect -406 32 -404 38
rect -397 32 -395 45
rect -308 58 -306 62
rect -298 58 -296 62
rect -257 60 -256 64
rect -193 62 -191 65
rect -183 62 -181 65
rect -257 58 -255 60
rect -248 58 -246 61
rect -369 32 -367 44
rect -342 31 -340 49
rect -332 31 -330 49
rect -220 57 -218 61
rect -257 44 -255 48
rect -406 0 -404 12
rect -397 9 -395 12
rect -369 8 -367 12
rect -468 -4 -466 0
rect -458 -4 -456 0
rect -308 20 -306 38
rect -298 20 -296 38
rect -257 35 -255 41
rect -248 35 -246 48
rect -159 61 -157 65
rect -149 61 -147 65
rect -220 35 -218 47
rect -193 34 -191 52
rect -183 34 -181 52
rect -257 3 -255 15
rect -248 12 -246 15
rect -220 11 -218 15
rect -308 -4 -306 0
rect -298 -4 -296 0
rect -159 23 -157 41
rect -149 23 -147 41
rect -159 -1 -157 3
rect -149 -1 -147 3
rect -193 -9 -191 -6
rect -183 -9 -181 -6
rect -502 -12 -500 -9
rect -492 -12 -490 -9
rect -342 -12 -340 -9
rect -332 -12 -330 -9
<< polycontact >>
rect -53 361 -49 365
rect -147 323 -143 327
rect -55 343 -51 347
rect -137 329 -133 333
rect -49 333 -45 337
rect -208 307 -204 311
rect -190 309 -186 313
rect -180 303 -176 307
rect -394 280 -390 284
rect -392 262 -388 266
rect -398 252 -394 256
rect -310 248 -306 252
rect -300 242 -296 246
rect -418 188 -414 192
rect -397 188 -393 192
rect -387 194 -383 198
rect -60 275 -56 279
rect -267 222 -263 226
rect -257 228 -253 232
rect -111 255 -107 259
rect -101 261 -97 265
rect -50 269 -46 273
rect -29 269 -25 273
rect -239 226 -235 230
rect -346 180 -342 184
rect -279 190 -275 194
rect -336 174 -332 178
rect -610 126 -606 130
rect -545 129 -541 133
rect -270 152 -266 156
rect -248 152 -244 156
rect -521 103 -517 107
rect -511 109 -507 113
rect -416 138 -412 142
rect -280 134 -276 138
rect -493 107 -489 111
rect -472 107 -468 111
rect -601 88 -597 92
rect -579 88 -575 92
rect -462 101 -458 105
rect -407 100 -403 104
rect -385 100 -381 104
rect -417 82 -413 86
rect -611 70 -607 74
rect -565 57 -561 61
rect -506 44 -502 48
rect -555 39 -551 43
rect -533 39 -529 43
rect -496 38 -492 42
rect -405 57 -401 61
rect -564 1 -560 5
rect -472 27 -468 31
rect -462 33 -458 37
rect -256 60 -252 64
rect -346 44 -342 48
rect -395 39 -391 43
rect -373 39 -369 43
rect -336 38 -332 42
rect -404 1 -400 5
rect -312 27 -308 31
rect -302 33 -298 37
rect -197 47 -193 51
rect -246 42 -242 46
rect -224 42 -220 46
rect -187 41 -183 45
rect -255 4 -251 8
rect -163 30 -159 34
rect -153 36 -149 40
<< metal1 >>
rect -90 376 -50 379
rect -206 367 -131 370
rect -90 370 -87 376
rect -53 372 -50 376
rect -118 367 -87 370
rect -60 369 -48 372
rect -206 349 -203 367
rect -178 360 -175 367
rect -154 360 -150 367
rect -135 360 -132 367
rect -230 346 -203 349
rect -393 295 -353 298
rect -393 291 -390 295
rect -395 288 -383 291
rect -356 289 -353 295
rect -356 286 -325 289
rect -230 289 -227 346
rect -206 338 -203 346
rect -145 339 -142 340
rect -154 336 -142 339
rect -154 327 -151 336
rect -118 333 -115 367
rect -133 330 -115 333
rect -107 360 -80 363
rect -112 335 -109 358
rect -53 354 -50 361
rect -38 360 -27 363
rect -30 354 -27 360
rect -62 351 -45 354
rect -48 345 -45 351
rect -34 351 -27 354
rect -112 332 -102 335
rect -172 324 -151 327
rect -215 311 -212 318
rect -197 311 -194 320
rect -172 313 -169 324
rect -154 322 -151 324
rect -143 323 -124 326
rect -127 320 -124 323
rect -112 322 -109 332
rect -55 326 -52 343
rect -48 342 -44 345
rect -30 336 -27 351
rect -49 331 -45 333
rect -34 332 -30 335
rect -49 329 -48 331
rect -112 319 -64 322
rect -222 308 -212 311
rect -215 306 -212 308
rect -204 308 -194 311
rect -186 310 -169 313
rect -112 312 -109 319
rect -67 316 -64 319
rect -67 313 -27 316
rect -197 306 -194 308
rect -197 303 -185 306
rect -176 304 -172 307
rect -188 302 -185 303
rect -61 306 -58 313
rect -43 306 -39 313
rect -135 297 -132 302
rect -30 300 -27 313
rect -312 286 -227 289
rect -206 288 -203 296
rect -197 288 -194 292
rect -178 288 -175 292
rect -171 294 -123 297
rect -171 288 -168 294
rect -416 279 -405 282
rect -416 273 -413 279
rect -393 273 -390 280
rect -363 279 -336 282
rect -416 270 -409 273
rect -416 255 -413 270
rect -398 270 -381 273
rect -398 264 -395 270
rect -399 261 -395 264
rect -413 251 -409 254
rect -397 247 -394 252
rect -445 243 -394 247
rect -391 245 -388 262
rect -334 254 -331 277
rect -341 251 -331 254
rect -334 241 -331 251
rect -328 252 -325 286
rect -311 279 -308 286
rect -293 279 -289 286
rect -268 279 -265 286
rect -301 258 -298 259
rect -301 255 -289 258
rect -328 249 -310 252
rect -292 246 -289 255
rect -240 257 -237 286
rect -215 285 -168 288
rect -379 238 -331 241
rect -314 242 -300 245
rect -292 243 -271 246
rect -292 241 -289 243
rect -379 235 -376 238
rect -455 232 -376 235
rect -562 169 -491 170
rect -562 167 -479 169
rect -562 166 -552 167
rect -562 139 -558 166
rect -546 160 -543 167
rect -522 160 -519 167
rect -494 166 -479 167
rect -494 148 -491 166
rect -482 159 -479 166
rect -455 159 -452 232
rect -416 219 -413 232
rect -404 225 -400 232
rect -385 225 -382 232
rect -334 231 -331 238
rect -274 232 -271 243
rect -274 229 -257 232
rect -249 230 -246 239
rect -231 230 -228 237
rect -249 227 -239 230
rect -271 223 -267 226
rect -249 225 -246 227
rect -231 227 -225 230
rect -231 225 -228 227
rect -258 222 -246 225
rect -258 221 -255 222
rect -311 216 -308 221
rect -320 213 -272 216
rect -395 204 -392 205
rect -404 201 -392 204
rect -425 192 -422 199
rect -404 192 -401 201
rect -383 195 -356 198
rect -428 189 -422 192
rect -425 187 -422 189
rect -414 189 -401 192
rect -404 187 -401 189
rect -393 188 -379 191
rect -359 182 -356 195
rect -353 182 -350 191
rect -359 179 -350 182
rect -342 181 -329 184
rect -416 163 -413 177
rect -353 177 -350 179
rect -353 174 -341 177
rect -332 175 -324 178
rect -344 173 -341 174
rect -419 160 -417 163
rect -482 156 -452 159
rect -385 162 -382 167
rect -412 159 -376 162
rect -353 159 -350 163
rect -334 159 -331 163
rect -320 159 -317 213
rect -275 207 -272 213
rect -268 207 -265 211
rect -249 207 -246 211
rect -240 207 -237 215
rect -215 207 -212 285
rect -126 240 -123 294
rect -51 285 -48 286
rect -51 282 -39 285
rect -87 276 -60 279
rect -114 262 -101 265
rect -93 263 -90 272
rect -87 263 -84 276
rect -42 273 -39 282
rect -21 273 -18 280
rect -74 269 -50 272
rect -42 270 -29 273
rect -74 267 -70 269
rect -42 268 -39 270
rect -21 270 -15 273
rect -21 268 -18 270
rect -93 260 -84 263
rect -120 258 -111 259
rect -115 256 -111 258
rect -93 258 -90 260
rect -102 255 -90 258
rect -102 254 -99 255
rect -112 240 -109 244
rect -93 240 -90 244
rect -61 243 -58 248
rect -30 244 -27 258
rect -67 240 -31 243
rect -126 237 -63 240
rect -275 204 -212 207
rect -275 191 -264 193
rect -275 190 -260 191
rect -263 183 -260 190
rect -249 183 -245 192
rect -265 180 -252 183
rect -380 156 -317 159
rect -285 156 -282 163
rect -277 162 -274 165
rect -450 148 -382 151
rect -494 145 -445 148
rect -635 135 -558 139
rect -635 62 -631 135
rect -606 126 -591 129
rect -594 119 -591 126
rect -580 119 -576 135
rect -537 133 -534 140
rect -494 138 -491 145
rect -473 138 -470 145
rect -455 138 -451 145
rect -386 143 -382 148
rect -400 141 -397 143
rect -412 138 -397 141
rect -400 135 -397 138
rect -386 140 -367 143
rect -549 130 -545 133
rect -537 130 -526 133
rect -400 131 -399 135
rect -537 128 -534 130
rect -596 116 -583 119
rect -616 92 -613 99
rect -608 98 -605 101
rect -625 90 -613 92
rect -620 89 -613 90
rect -616 86 -613 89
rect -608 86 -605 93
rect -586 92 -583 116
rect -597 88 -594 91
rect -586 89 -579 92
rect -596 75 -590 79
rect -596 73 -595 75
rect -607 70 -595 73
rect -635 58 -593 62
rect -586 61 -583 89
rect -571 83 -568 99
rect -571 81 -567 83
rect -568 78 -567 81
rect -580 72 -577 77
rect -546 72 -543 118
rect -529 113 -526 130
rect -402 130 -399 131
rect -386 131 -382 140
rect -394 130 -389 131
rect -402 128 -389 130
rect -529 110 -511 113
rect -503 111 -500 120
rect -485 111 -482 118
rect -463 117 -460 118
rect -463 114 -451 117
rect -503 108 -493 111
rect -524 104 -521 107
rect -503 106 -500 108
rect -485 108 -472 111
rect -485 106 -482 108
rect -512 103 -500 106
rect -512 102 -509 103
rect -454 105 -451 114
rect -474 101 -462 104
rect -454 104 -431 105
rect -422 104 -419 111
rect -414 110 -411 113
rect -454 102 -419 104
rect -454 100 -451 102
rect -522 88 -519 92
rect -503 88 -500 92
rect -494 89 -491 96
rect -447 92 -444 102
rect -434 101 -431 102
rect -426 101 -419 102
rect -422 98 -419 101
rect -414 98 -411 105
rect -392 104 -389 128
rect -403 100 -400 103
rect -392 101 -385 104
rect -377 95 -374 111
rect -377 93 -373 95
rect -533 85 -495 88
rect -533 72 -530 85
rect -402 87 -396 91
rect -402 85 -401 87
rect -413 82 -401 85
rect -374 90 -373 93
rect -386 84 -383 89
rect -364 84 -361 156
rect -297 154 -282 156
rect -297 153 -294 154
rect -289 153 -282 154
rect -285 150 -282 153
rect -277 150 -274 157
rect -255 156 -252 180
rect -266 152 -263 155
rect -255 153 -248 156
rect -240 147 -237 163
rect -240 145 -236 147
rect -265 139 -259 143
rect -265 137 -264 139
rect -276 134 -264 137
rect -237 142 -236 145
rect -249 136 -246 141
rect -249 133 -244 136
rect -249 129 -246 133
rect -334 126 -246 129
rect -334 94 -331 126
rect -334 91 -268 94
rect -386 81 -361 84
rect -473 76 -470 80
rect -580 69 -530 72
rect -364 75 -361 81
rect -271 79 -268 91
rect -469 72 -361 75
rect -534 66 -530 69
rect -364 66 -361 72
rect -294 76 -222 79
rect -294 66 -291 76
rect -534 63 -470 66
rect -597 -15 -593 58
rect -561 58 -549 61
rect -550 56 -549 58
rect -550 52 -544 56
rect -534 54 -531 63
rect -507 59 -504 63
rect -488 59 -485 63
rect -524 54 -521 56
rect -522 50 -521 54
rect -473 58 -470 63
rect -374 63 -291 66
rect -225 69 -222 76
rect -225 66 -142 69
rect -401 58 -389 61
rect -390 56 -389 58
rect -582 41 -579 42
rect -570 42 -567 45
rect -574 41 -567 42
rect -582 39 -567 41
rect -582 -4 -579 39
rect -570 32 -567 39
rect -562 38 -559 45
rect -551 40 -548 43
rect -540 39 -533 42
rect -540 35 -537 39
rect -562 30 -559 33
rect -525 32 -522 50
rect -390 52 -384 56
rect -374 54 -371 63
rect -347 59 -344 63
rect -328 59 -325 63
rect -364 54 -361 56
rect -362 50 -361 54
rect -313 58 -310 63
rect -497 48 -494 49
rect -509 44 -506 47
rect -497 47 -485 48
rect -497 45 -482 47
rect -488 44 -477 45
rect -513 38 -496 41
rect -513 35 -510 38
rect -540 15 -537 30
rect -488 31 -485 44
rect -475 34 -462 37
rect -454 36 -451 38
rect -422 41 -419 42
rect -410 42 -407 45
rect -414 41 -407 42
rect -422 39 -407 41
rect -448 36 -445 39
rect -454 33 -445 36
rect -479 27 -472 30
rect -479 23 -476 27
rect -454 24 -451 33
rect -463 21 -451 24
rect -463 20 -460 21
rect -550 12 -537 15
rect -548 5 -545 12
rect -560 2 -545 5
rect -534 3 -530 12
rect -549 -4 -546 2
rect -534 0 -510 3
rect -513 -15 -510 0
rect -597 -16 -510 -15
rect -473 -7 -470 0
rect -455 -7 -451 0
rect -422 -4 -419 39
rect -410 32 -407 39
rect -402 38 -399 45
rect -391 40 -388 43
rect -380 39 -373 42
rect -380 35 -377 39
rect -402 30 -399 33
rect -365 32 -362 50
rect -337 48 -334 49
rect -349 44 -346 47
rect -337 47 -325 48
rect -337 45 -322 47
rect -328 44 -317 45
rect -353 38 -336 41
rect -353 35 -350 38
rect -380 15 -377 30
rect -328 31 -325 44
rect -315 34 -302 37
rect -294 36 -291 38
rect -288 36 -285 66
rect -252 61 -240 64
rect -241 59 -240 61
rect -241 55 -235 59
rect -225 57 -222 66
rect -198 62 -195 66
rect -179 62 -176 66
rect -215 57 -212 59
rect -213 53 -212 57
rect -164 61 -161 66
rect -294 33 -285 36
rect -273 44 -270 45
rect -261 45 -258 48
rect -265 44 -258 45
rect -273 42 -258 44
rect -319 27 -312 30
rect -319 23 -316 27
rect -294 24 -291 33
rect -303 21 -291 24
rect -303 20 -300 21
rect -390 12 -377 15
rect -388 5 -385 12
rect -400 2 -385 5
rect -374 3 -370 12
rect -389 -4 -386 2
rect -374 0 -350 3
rect -507 -16 -504 -9
rect -483 -10 -445 -7
rect -483 -15 -479 -10
rect -353 -15 -350 0
rect -483 -16 -350 -15
rect -313 -7 -310 0
rect -295 -7 -291 0
rect -273 -1 -270 42
rect -261 35 -258 42
rect -253 41 -250 48
rect -242 43 -239 46
rect -231 42 -224 45
rect -231 38 -228 42
rect -253 33 -250 36
rect -216 35 -213 53
rect -188 51 -185 52
rect -200 47 -197 50
rect -188 50 -176 51
rect -188 48 -173 50
rect -179 47 -168 48
rect -204 41 -187 44
rect -204 38 -201 41
rect -231 18 -228 33
rect -179 34 -176 47
rect -166 37 -153 40
rect -145 39 -142 41
rect -139 39 -136 76
rect -145 36 -136 39
rect -170 30 -163 33
rect -170 26 -167 30
rect -145 27 -142 36
rect -154 24 -142 27
rect -154 23 -151 24
rect -241 15 -228 18
rect -239 8 -236 15
rect -251 5 -236 8
rect -225 6 -221 15
rect -240 -1 -237 5
rect -225 3 -201 6
rect -204 -7 -201 3
rect -347 -16 -344 -9
rect -323 -10 -201 -7
rect -323 -16 -319 -10
rect -204 -13 -201 -10
rect -164 -4 -161 3
rect -146 -4 -142 3
rect -198 -13 -195 -6
rect -174 -7 -136 -4
rect -174 -13 -170 -7
rect -204 -16 -170 -13
rect -597 -19 -319 -16
<< m2contact >>
rect -131 367 -126 372
rect -317 286 -312 291
rect -112 358 -107 363
rect -128 315 -123 320
rect -57 321 -52 326
rect -336 277 -331 282
rect -391 240 -386 245
rect -225 226 -220 231
rect -433 187 -428 192
rect -329 181 -324 186
rect -15 268 -10 273
rect -264 191 -259 196
rect -278 157 -273 162
rect -609 93 -604 98
rect -595 70 -590 75
rect -567 78 -562 83
rect -399 130 -394 135
rect -415 105 -410 110
rect -495 84 -490 89
rect -401 82 -396 87
rect -373 90 -368 95
rect -264 134 -259 139
rect -236 142 -231 147
rect -474 71 -469 76
rect -140 76 -135 81
rect -587 56 -582 61
rect -549 56 -544 61
rect -521 53 -516 58
rect -288 66 -283 72
rect -389 56 -384 61
rect -563 33 -558 38
rect -541 30 -536 35
rect -361 53 -356 58
rect -482 45 -477 50
rect -514 30 -509 35
rect -480 33 -475 38
rect -403 33 -398 38
rect -381 30 -376 35
rect -322 45 -317 50
rect -354 30 -349 35
rect -320 33 -315 38
rect -240 59 -235 64
rect -212 56 -207 61
rect -254 36 -249 41
rect -232 33 -227 38
rect -205 33 -200 38
rect -171 36 -166 41
<< metal2 >>
rect -628 97 -625 578
rect -441 109 -438 576
rect -126 368 -109 371
rect -112 363 -109 368
rect -119 322 -57 325
rect -334 287 -317 290
rect -334 282 -331 287
rect -126 284 -123 315
rect -245 279 -234 282
rect -245 262 -242 279
rect -210 281 -123 284
rect -327 259 -242 262
rect -327 244 -324 259
rect -386 241 -324 244
rect -432 226 -373 229
rect -432 192 -429 226
rect -327 186 -324 241
rect -318 191 -315 240
rect -224 199 -221 226
rect -263 196 -221 199
rect -318 188 -305 191
rect -324 181 -313 184
rect -316 155 -313 181
rect -359 152 -313 155
rect -400 130 -399 133
rect -394 130 -390 133
rect -393 126 -390 130
rect -441 106 -415 109
rect -628 94 -609 97
rect -593 68 -590 70
rect -566 68 -563 78
rect -593 65 -563 68
rect -529 68 -526 102
rect -490 85 -474 88
rect -477 72 -474 85
rect -399 80 -396 82
rect -372 80 -369 90
rect -399 77 -369 80
rect -359 71 -356 152
rect -308 148 -305 188
rect -300 161 -296 194
rect -210 190 -207 281
rect -119 267 -116 322
rect -70 307 -11 310
rect -14 273 -11 307
rect -227 187 -207 190
rect -300 158 -278 161
rect -352 145 -305 148
rect -352 79 -349 145
rect -293 139 -290 149
rect -342 136 -290 139
rect -342 87 -339 136
rect -262 132 -259 134
rect -235 132 -232 142
rect -262 129 -232 132
rect -227 124 -224 187
rect -328 121 -224 124
rect -328 99 -325 121
rect -328 96 -263 99
rect -342 84 -274 87
rect -352 76 -284 79
rect -287 72 -284 76
rect -359 68 -318 71
rect -529 65 -478 68
rect -544 56 -521 57
rect -586 37 -583 56
rect -548 54 -521 56
rect -481 50 -478 65
rect -586 34 -563 37
rect -513 37 -510 39
rect -513 35 -480 37
rect -536 31 -514 34
rect -509 34 -480 35
rect -426 37 -423 57
rect -384 56 -361 57
rect -388 54 -361 56
rect -321 50 -318 68
rect -277 40 -274 84
rect -266 84 -263 96
rect -266 81 -215 84
rect -218 80 -215 81
rect -218 77 -140 80
rect -235 59 -212 60
rect -239 57 -212 59
rect -426 34 -403 37
rect -353 37 -350 39
rect -353 35 -320 37
rect -376 31 -354 34
rect -349 34 -320 35
rect -277 37 -254 40
rect -204 40 -201 42
rect -204 38 -171 40
rect -227 34 -205 37
rect -200 37 -171 38
<< m3contact >>
rect -373 225 -368 230
rect -75 306 -70 311
<< m123contact >>
rect -450 242 -445 247
rect -554 129 -549 134
rect -30 331 -25 336
rect -48 326 -43 331
rect -172 302 -167 307
rect -418 250 -413 255
rect -379 186 -374 191
rect -319 240 -314 245
rect -276 221 -271 226
rect -328 170 -323 175
rect -417 158 -412 163
rect -529 102 -524 107
rect -625 85 -620 90
rect -594 87 -589 92
rect -479 99 -474 104
rect -431 97 -426 102
rect -400 99 -395 104
rect -448 87 -443 92
rect -119 262 -114 267
rect -75 262 -70 267
rect -120 253 -115 258
rect -31 239 -26 244
rect -294 149 -289 154
rect -263 151 -258 156
rect -579 41 -574 46
rect -514 44 -509 49
rect -548 39 -543 44
rect -448 39 -443 44
rect -419 41 -414 46
rect -354 44 -349 49
rect -388 39 -383 44
rect -270 44 -265 49
rect -205 47 -200 52
rect -173 48 -168 53
rect -239 42 -234 47
rect -480 18 -475 23
rect -320 18 -315 23
rect -171 21 -166 26
<< metal3 >>
rect -237 326 -48 329
rect -237 297 -234 326
rect -76 311 -69 312
rect -76 310 -75 311
rect -168 307 -75 310
rect -167 304 -165 307
rect -76 306 -75 307
rect -70 306 -69 311
rect -76 305 -69 306
rect -318 294 -234 297
rect -553 182 -498 185
rect -553 134 -550 182
rect -501 181 -498 182
rect -501 178 -477 181
rect -529 173 -513 176
rect -593 130 -554 133
rect -593 92 -590 130
rect -529 107 -526 173
rect -448 154 -445 242
rect -417 163 -414 250
rect -318 245 -315 294
rect -204 275 -129 278
rect -374 230 -367 231
rect -374 225 -373 230
rect -368 229 -367 230
rect -368 226 -275 229
rect -368 225 -367 226
rect -374 224 -367 225
rect -278 223 -276 226
rect -374 186 -372 191
rect -375 173 -372 186
rect -204 183 -201 275
rect -132 266 -129 275
rect -132 263 -119 266
rect -136 255 -120 258
rect -74 236 -71 262
rect -29 244 -26 331
rect -138 233 -71 236
rect -221 180 -201 183
rect -375 170 -364 173
rect -372 169 -369 170
rect -478 151 -445 154
rect -478 104 -475 151
rect -328 153 -324 170
rect -292 154 -263 155
rect -400 149 -324 153
rect -289 152 -263 154
rect -221 118 -218 180
rect -320 115 -218 118
rect -320 105 -317 115
rect -429 102 -400 103
rect -623 90 -594 91
rect -620 88 -594 90
rect -551 44 -514 47
rect -478 44 -475 99
rect -426 100 -400 102
rect -320 102 -256 105
rect -259 92 -256 102
rect -443 87 -439 91
rect -259 89 -208 92
rect -442 86 -439 87
rect -211 86 -208 89
rect -442 83 -441 86
rect -211 83 -169 86
rect -172 53 -169 83
rect -551 43 -548 44
rect -574 41 -548 43
rect -577 40 -548 41
rect -513 22 -510 44
rect -478 41 -448 44
rect -391 44 -354 47
rect -242 47 -205 50
rect -242 46 -239 47
rect -265 44 -239 46
rect -391 43 -388 44
rect -414 41 -388 43
rect -417 40 -388 41
rect -513 19 -480 22
rect -353 22 -350 44
rect -268 43 -239 44
rect -204 25 -201 47
rect -353 19 -320 22
rect -204 22 -171 25
<< m234contact >>
rect -234 278 -229 283
rect -301 194 -296 199
rect -405 149 -400 154
rect -394 121 -389 126
rect -427 57 -422 62
<< m4contact >>
rect -477 177 -472 182
rect -513 172 -508 177
rect -141 255 -136 260
rect -369 165 -364 170
<< metal4 >>
rect -300 199 -297 296
rect -229 278 -224 282
rect -227 272 -224 278
rect -227 269 -141 272
rect -144 255 -141 269
rect -472 179 -376 182
rect -508 173 -484 176
rect -487 153 -484 173
rect -379 168 -376 179
rect -379 165 -369 168
rect -487 150 -405 153
rect -393 70 -390 121
rect -426 67 -390 70
rect -426 62 -423 67
<< m345contact >>
rect -143 232 -138 237
rect -441 81 -436 86
<< metal5 >>
rect -198 264 -146 267
rect -198 193 -195 264
rect -149 237 -146 264
rect -149 233 -143 237
rect -225 190 -195 193
rect -225 147 -222 190
rect -357 144 -222 147
rect -357 85 -354 144
rect -436 82 -354 85
<< labels >>
rlabel metal1 -554 60 -554 60 1 b0_inv
rlabel metal1 -451 33 -445 36 7 g0_inv
rlabel metal1 -485 44 -481 47 1 p0_inv
rlabel metal1 -548 -2 -546 1 1 b0
rlabel metal2 -586 58 -584 60 3 mid_s0
rlabel metal1 -573 39 -571 41 1 a0
rlabel metal1 -506 -18 -506 -17 1 vdd
rlabel metal1 -496 64 -496 64 5 gnd
rlabel metal1 -576 70 -576 70 1 gnd
rlabel metal1 -607 91 -605 93 1 s0
rlabel metal1 -619 90 -617 92 1 c0
rlabel metal1 -586 89 -583 91 1 mid_s0
rlabel metal1 -451 102 -445 105 7 c1
rlabel metal1 -478 102 -474 104 1 g0_inv
rlabel metal1 -458 73 -458 73 1 gnd
rlabel metal1 -484 109 -482 112 1 temp100
rlabel metal1 -511 87 -511 87 1 gnd
rlabel metal1 -536 131 -534 134 1 c0_inv
rlabel metal1 -551 130 -549 132 3 c0
rlabel metal1 -361 2 -361 2 1 vdd
rlabel metal1 -336 64 -336 64 5 gnd
rlabel metal1 -346 -18 -346 -17 1 vdd
rlabel metal1 -307 -8 -307 -8 1 vdd
rlabel metal2 -426 58 -424 60 3 mid_s1
rlabel metal1 -413 39 -411 41 1 a1
rlabel metal1 -388 -2 -386 1 1 b1
rlabel metal1 -325 44 -321 47 1 p1_inv
rlabel metal1 -291 33 -285 36 7 g1_inv
rlabel m2contact -387 59 -385 61 1 b1_inv
rlabel metal1 -413 103 -411 105 1 s1
rlabel metal1 -373 141 -373 141 5 vdd
rlabel metal1 -332 239 -332 240 5 vdd
rlabel metal1 -342 158 -342 158 1 gnd
rlabel metal1 -331 181 -327 183 7 p1_inv
rlabel metal1 -330 175 -325 177 7 p0_inv
rlabel metal1 -358 179 -354 181 3 temp101
rlabel metal1 -388 233 -388 233 5 vdd
rlabel metal1 -397 160 -397 160 1 gnd
rlabel metal1 -381 189 -377 190 1 c0
rlabel metal1 -425 190 -423 192 1 temp102
rlabel metal1 -414 262 -414 262 3 gnd
rlabel metal1 -333 252 -332 252 7 vdd
rlabel metal1 -392 288 -389 291 1 temp103
rlabel metal1 -305 287 -305 287 5 vdd
rlabel metal1 -296 214 -296 214 1 gnd
rlabel metal1 -313 243 -313 243 1 g1_inv
rlabel metal1 -289 243 -283 246 7 temp104
rlabel metal1 -267 287 -267 288 5 vdd
rlabel metal1 -257 206 -257 206 1 gnd
rlabel metal1 -230 228 -228 230 1 c2
rlabel metal1 -397 244 -394 247 1 g0_inv
rlabel metal1 -528 104 -523 107 1 p0_inv
rlabel metal1 -239 1 -237 4 1 b2
rlabel metal1 -264 42 -262 44 1 a2
rlabel metal2 -277 61 -275 63 3 mid_s2
rlabel m2contact -238 62 -236 64 1 b2_inv
rlabel metal1 -176 47 -172 50 1 p2_inv
rlabel metal1 -142 36 -136 39 7 g2_inv
rlabel metal1 -158 -5 -158 -5 1 vdd
rlabel metal1 -197 -15 -197 -14 1 vdd
rlabel metal1 -187 67 -187 67 5 gnd
rlabel metal1 -212 5 -212 5 1 vdd
rlabel metal1 -276 155 -274 157 1 s2
rlabel metal1 -245 134 -245 134 1 gnd
rlabel metal1 -111 320 -111 321 5 vdd
rlabel metal1 -101 239 -101 239 1 gnd
rlabel metal1 -55 314 -55 314 5 vdd
rlabel metal1 -46 241 -46 241 1 gnd
rlabel metal1 -29 343 -29 343 7 gnd
rlabel metal1 -111 333 -110 333 3 vdd
rlabel metal1 -138 368 -138 368 5 vdd
rlabel metal1 -147 295 -147 295 1 gnd
rlabel metal1 -176 368 -176 369 5 vdd
rlabel metal1 -186 287 -186 287 1 gnd
rlabel metal1 -215 309 -213 311 1 c3
rlabel metal1 -160 324 -154 327 1 temp108
rlabel metal1 -20 271 -18 273 1 temp106
rlabel metal1 -66 270 -62 271 1 c1
rlabel metal1 -89 260 -85 262 1 temp105
rlabel metal1 -116 262 -112 264 1 p2_inv
rlabel metal1 -54 369 -51 372 1 temp107
rlabel metal1 -131 323 -129 325 1 g2_inv
rlabel metal1 -48 327 -45 330 1 g1_inv
rlabel metal1 -114 257 -114 257 1 p1_inv
<< end >>
