* SPICE3 file created from XOR.ext - technology: scmos

.option scale=0.09u

M1000 vdd in1 in1_inv w_n60_18# pfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 in2 in1 out w_n21_23# pfet w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1002 out in2 in1 w_n21_23# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1003 gnd in1 in1_inv Gnd nfet w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1004 out in2 in1_inv Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1005 in2 in1_inv out Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 w_n60_18# in1_inv 0.02fF
C1 w_n21_23# in1 0.10fF
C2 in1 in1_inv 0.06fF
C3 in1 in2 0.03fF
C4 w_n21_23# out 0.17fF
C5 w_n60_18# vdd 0.02fF
C6 w_n60_18# in1 0.07fF
C7 in2 out 0.34fF
C8 w_n21_23# in2 0.09fF
C9 in2 in1_inv 0.10fF
C10 in1 out 0.00fF
C11 in1 gnd 0.02fF
C12 out Gnd 0.07fF
C13 in1_inv Gnd 0.03fF
C14 vdd Gnd 0.01fF
C15 gnd Gnd 0.03fF
C16 in2 Gnd 0.41fF
C17 in1 Gnd 0.13fF
C18 w_n21_23# Gnd 0.53fF
C19 w_n60_18# Gnd 0.80fF
