magic
tech scmos
timestamp 1731409616
<< nwell >>
rect -176 109 -99 131
rect -59 125 -27 144
rect -194 99 -99 109
rect -81 119 -27 125
rect -194 79 -142 99
rect -81 91 -29 119
rect -194 77 -170 79
rect -91 31 -57 83
rect -40 71 -6 77
rect -40 45 16 71
rect -9 39 16 45
<< ntransistor >>
rect -21 130 -11 132
rect -17 112 -7 114
rect -17 102 -7 104
rect -183 61 -181 71
rect -122 67 -120 87
rect -112 67 -110 87
rect -165 57 -163 67
rect -155 57 -153 67
rect -80 9 -78 19
rect -70 9 -68 19
rect -29 13 -27 33
rect -19 13 -17 33
rect 2 23 4 33
<< ptransistor >>
rect -53 130 -33 132
rect -183 83 -181 103
rect -165 85 -163 125
rect -155 85 -153 125
rect -122 105 -120 125
rect -112 105 -110 125
rect -75 112 -35 114
rect -75 102 -35 104
rect -80 37 -78 77
rect -70 37 -68 77
rect -29 51 -27 71
rect -19 51 -17 71
rect 2 45 4 65
<< ndiffusion >>
rect -17 133 -11 137
rect -21 132 -11 133
rect -21 129 -11 130
rect -21 125 -15 129
rect -17 115 -11 119
rect -17 114 -7 115
rect -17 110 -7 112
rect -13 106 -7 110
rect -17 104 -7 106
rect -17 101 -7 102
rect -17 97 -11 101
rect -184 67 -183 71
rect -188 61 -183 67
rect -181 65 -176 71
rect -123 83 -122 87
rect -127 67 -122 83
rect -120 67 -112 87
rect -110 71 -105 87
rect -110 67 -109 71
rect -181 61 -180 65
rect -170 61 -165 67
rect -166 57 -165 61
rect -163 63 -161 67
rect -157 63 -155 67
rect -163 57 -155 63
rect -153 61 -148 67
rect -153 57 -152 61
rect -85 13 -80 19
rect -81 9 -80 13
rect -78 15 -76 19
rect -72 15 -70 19
rect -78 9 -70 15
rect -68 13 -63 19
rect -34 17 -29 33
rect -30 13 -29 17
rect -27 13 -19 33
rect -17 29 -16 33
rect -17 13 -12 29
rect -3 27 2 33
rect 1 23 2 27
rect 4 29 5 33
rect 4 23 9 29
rect -68 9 -67 13
<< pdiffusion >>
rect -53 133 -37 137
rect -53 132 -33 133
rect -53 129 -33 130
rect -49 125 -33 129
rect -188 87 -183 103
rect -184 83 -183 87
rect -181 99 -180 103
rect -181 83 -176 99
rect -170 89 -165 125
rect -166 85 -165 89
rect -163 85 -155 125
rect -153 121 -152 125
rect -153 85 -148 121
rect -123 121 -122 125
rect -127 105 -122 121
rect -120 109 -112 125
rect -120 105 -118 109
rect -114 105 -112 109
rect -110 121 -109 125
rect -110 105 -105 121
rect -75 115 -39 119
rect -75 114 -35 115
rect -75 104 -35 112
rect -75 101 -35 102
rect -71 97 -35 101
rect -81 73 -80 77
rect -85 37 -80 73
rect -78 37 -70 77
rect -68 41 -63 77
rect -30 67 -29 71
rect -34 51 -29 67
rect -27 55 -19 71
rect -27 51 -25 55
rect -21 51 -19 55
rect -17 67 -16 71
rect -17 51 -12 67
rect 1 61 2 65
rect -68 37 -67 41
rect -3 45 2 61
rect 4 49 9 65
rect 4 45 5 49
<< ndcontact >>
rect -21 133 -17 137
rect -15 125 -11 129
rect -11 115 -7 119
rect -17 106 -13 110
rect -11 97 -7 101
rect -188 67 -184 71
rect -127 83 -123 87
rect -109 67 -105 71
rect -180 61 -176 65
rect -170 57 -166 61
rect -161 63 -157 67
rect -152 57 -148 61
rect -85 9 -81 13
rect -76 15 -72 19
rect -34 13 -30 17
rect -16 29 -12 33
rect -3 23 1 27
rect 5 29 9 33
rect -67 9 -63 13
<< pdcontact >>
rect -37 133 -33 137
rect -53 125 -49 129
rect -188 83 -184 87
rect -180 99 -176 103
rect -170 85 -166 89
rect -152 121 -148 125
rect -127 121 -123 125
rect -118 105 -114 109
rect -109 121 -105 125
rect -39 115 -35 119
rect -75 97 -71 101
rect -85 73 -81 77
rect -34 67 -30 71
rect -25 51 -21 55
rect -16 67 -12 71
rect -3 61 1 65
rect -67 37 -63 41
rect 5 45 9 49
<< polysilicon >>
rect -56 130 -53 132
rect -33 130 -21 132
rect -11 130 -8 132
rect -165 125 -163 128
rect -155 125 -153 128
rect -122 125 -120 129
rect -112 125 -110 129
rect -183 103 -181 106
rect -78 112 -75 114
rect -35 112 -17 114
rect -7 112 -4 114
rect -122 87 -120 105
rect -112 87 -110 105
rect -78 102 -75 104
rect -35 102 -17 104
rect -7 102 -4 104
rect -183 71 -181 83
rect -165 67 -163 85
rect -155 67 -153 85
rect -80 77 -78 80
rect -70 77 -68 80
rect -183 58 -181 61
rect -122 63 -120 67
rect -112 63 -110 67
rect -165 54 -163 57
rect -155 54 -153 57
rect -29 71 -27 75
rect -19 71 -17 75
rect 2 65 4 69
rect -80 19 -78 37
rect -70 19 -68 37
rect -29 33 -27 51
rect -19 33 -17 51
rect 2 33 4 45
rect 2 19 4 23
rect -29 9 -27 13
rect -19 9 -17 13
rect -80 6 -78 9
rect -70 6 -68 9
<< polycontact >>
rect -26 126 -22 130
rect -120 88 -116 92
rect -28 108 -24 112
rect -110 94 -106 98
rect -22 98 -18 102
rect -181 72 -177 76
rect -163 74 -159 78
rect -153 68 -149 72
rect -33 40 -29 44
rect -84 20 -80 24
rect -74 26 -70 30
rect -23 34 -19 38
rect -2 34 2 38
<< metal1 >>
rect -63 141 -23 144
rect -179 132 -104 135
rect -63 135 -60 141
rect -26 137 -23 141
rect -91 132 -60 135
rect -33 134 -21 137
rect -179 103 -176 132
rect -151 125 -148 132
rect -127 125 -123 132
rect -108 125 -105 132
rect -118 104 -115 105
rect -127 101 -115 104
rect -127 92 -124 101
rect -91 98 -88 132
rect -106 95 -88 98
rect -80 125 -53 128
rect -85 100 -82 123
rect -26 119 -23 126
rect -11 125 0 128
rect -3 119 0 125
rect -35 116 -18 119
rect -21 110 -18 116
rect -7 116 0 119
rect -85 97 -75 100
rect -145 89 -124 92
rect -188 76 -185 83
rect -170 76 -167 85
rect -145 78 -142 89
rect -127 87 -124 89
rect -116 88 -99 91
rect -85 87 -82 97
rect -28 91 -25 108
rect -21 107 -17 110
rect -3 101 0 116
rect -22 91 -19 98
rect -7 97 -3 100
rect -85 84 -37 87
rect -195 73 -185 76
rect -188 71 -185 73
rect -177 73 -167 76
rect -159 75 -142 78
rect -85 77 -82 84
rect -40 81 -37 84
rect -40 78 0 81
rect -170 71 -167 73
rect -170 68 -158 71
rect -149 69 -145 72
rect -161 67 -158 68
rect -34 71 -31 78
rect -16 71 -12 78
rect -108 62 -105 67
rect -3 65 0 78
rect -179 53 -176 61
rect -170 53 -167 57
rect -151 53 -148 57
rect -144 59 -96 62
rect -144 53 -141 59
rect -179 50 -141 53
rect -99 5 -96 59
rect -24 50 -21 51
rect -24 47 -12 50
rect -60 41 -33 44
rect -87 27 -74 30
rect -66 28 -63 37
rect -60 28 -57 41
rect -15 38 -12 47
rect 6 38 9 45
rect -40 34 -23 37
rect -15 35 -2 38
rect -15 33 -12 35
rect 6 35 12 38
rect 6 33 9 35
rect -66 25 -57 28
rect -92 21 -84 24
rect -66 23 -63 25
rect -75 20 -63 23
rect -75 19 -72 20
rect -85 5 -82 9
rect -66 5 -63 9
rect -34 8 -31 13
rect -3 9 0 23
rect -40 5 -4 8
rect -99 2 -36 5
<< m2contact >>
rect -104 132 -99 137
rect -85 123 -80 128
rect -30 86 -25 91
rect -92 27 -87 32
rect 12 33 17 38
rect -93 16 -88 21
<< metal2 >>
rect -99 133 -82 136
rect -85 128 -82 133
rect -92 87 -30 90
rect -92 32 -89 87
rect -43 72 16 75
rect 13 38 16 72
<< m3contact >>
rect -48 71 -43 76
<< m123contact >>
rect -3 96 2 101
rect -145 67 -140 72
rect -4 4 1 9
<< metal3 >>
rect -49 76 -42 77
rect -49 75 -48 76
rect -141 72 -48 75
rect -140 69 -138 72
rect -49 71 -48 72
rect -43 71 -42 76
rect -49 70 -42 71
rect -2 9 1 96
<< labels >>
rlabel metal1 -84 85 -84 86 5 vdd
rlabel metal1 -74 4 -74 4 1 gnd
rlabel metal1 -89 27 -85 29 3 p1_inv
rlabel metal1 -91 21 -86 23 3 p0_inv
rlabel metal1 -62 25 -58 27 7 temp101
rlabel metal1 -28 79 -28 79 5 vdd
rlabel metal1 -19 6 -19 6 1 gnd
rlabel metal1 -39 35 -35 36 1 c0
rlabel metal1 7 36 9 38 1 temp102
rlabel metal1 -2 108 -2 108 7 gnd
rlabel metal1 -84 98 -83 98 3 vdd
rlabel metal1 -22 92 -19 95 1 g0_inv
rlabel metal1 -27 134 -24 137 1 temp103
rlabel metal1 -111 133 -111 133 5 vdd
rlabel metal1 -120 60 -120 60 1 gnd
rlabel metal1 -103 89 -103 89 1 g1_inv
rlabel metal1 -133 89 -127 92 3 temp104
rlabel metal1 -149 133 -149 134 5 vdd
rlabel metal1 -159 52 -159 52 1 gnd
rlabel metal1 -188 74 -186 76 1 c2
<< end >>
