magic
tech scmos
timestamp 1731426413
<< nwell >>
rect -67 39 1 71
<< ntransistor >>
rect -56 7 -54 27
rect -46 7 -44 27
rect -22 7 -20 27
rect -12 7 -10 27
<< ptransistor >>
rect -56 45 -54 65
rect -46 45 -44 65
rect -22 45 -20 65
rect -12 45 -10 65
<< ndiffusion >>
rect -61 11 -56 27
rect -57 7 -56 11
rect -54 7 -46 27
rect -44 23 -43 27
rect -44 7 -39 23
rect -27 11 -22 27
rect -23 7 -22 11
rect -20 7 -12 27
rect -10 23 -9 27
rect -10 7 -5 23
<< pdiffusion >>
rect -57 61 -56 65
rect -61 45 -56 61
rect -54 49 -46 65
rect -54 45 -52 49
rect -48 45 -46 49
rect -44 61 -43 65
rect -44 45 -39 61
rect -23 61 -22 65
rect -27 45 -22 61
rect -20 49 -12 65
rect -20 45 -18 49
rect -14 45 -12 49
rect -10 61 -9 65
rect -10 45 -5 61
<< ndcontact >>
rect -61 7 -57 11
rect -43 23 -39 27
rect -27 7 -23 11
rect -9 23 -5 27
<< pdcontact >>
rect -61 61 -57 65
rect -52 45 -48 49
rect -43 61 -39 65
rect -27 61 -23 65
rect -18 45 -14 49
rect -9 61 -5 65
<< polysilicon >>
rect -56 65 -54 69
rect -46 65 -44 69
rect -22 65 -20 69
rect -12 65 -10 69
rect -56 27 -54 45
rect -46 27 -44 45
rect -22 27 -20 45
rect -12 27 -10 45
rect -56 3 -54 7
rect -46 3 -44 7
rect -22 3 -20 7
rect -12 3 -10 7
<< polycontact >>
rect -60 34 -56 38
rect -50 28 -46 32
rect -26 34 -22 38
rect -16 28 -12 32
<< metal1 >>
rect -67 72 1 75
rect -61 65 -58 72
rect -43 65 -39 72
rect -27 65 -24 72
rect -9 65 -5 72
rect -51 44 -48 45
rect -17 44 -14 45
rect -51 41 -39 44
rect -17 41 -5 44
rect -67 35 -60 38
rect -67 28 -50 31
rect -42 31 -39 41
rect -28 34 -26 38
rect -8 32 -5 41
rect -42 28 -16 31
rect -8 29 1 32
rect -42 27 -39 28
rect -8 27 -5 29
rect -61 2 -58 7
rect -27 2 -24 7
rect -67 -1 -2 2
<< m2contact >>
rect -33 34 -28 39
<< labels >>
rlabel metal1 -55 73 -55 73 5 vdd
rlabel metal1 -46 0 -46 0 1 gnd
rlabel metal1 -64 35 -62 38 3 p4
rlabel metal1 -65 28 -62 31 3 c0
rlabel metal1 -21 73 -21 73 5 vdd
rlabel metal1 -12 0 -12 0 1 gnd
rlabel metal1 -29 29 -27 30 1 temp113
rlabel m2contact -31 35 -28 38 1 g4_inv
rlabel metal1 -5 29 1 32 7 c4
<< end >>
