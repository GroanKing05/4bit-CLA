* SPICE3 file created from ThreeBitAdder.ext - technology: scmos

.option scale=0.09u

M1000 s0 c0 mid_s0 w_186_n314# pfet w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1001 mid_s0 a_41_n338# a0 Gnd nfet w=10 l=2
+  ad=70 pd=34 as=50 ps=30
M1002 a_636_n229# b2 vdd w_589_n235# pfet w=40 l=2
+  ad=320 pd=96 as=5120 ps=2412
M1003 p2_inv b2 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=2500 ps=1420
M1004 vdd mid_s2 a_632_n320# w_648_n327# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1005 gnd temp101 a_410_n252# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1006 gnd a_387_n246# temp102 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1007 gnd temp107 a_744_n230# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1008 a_546_n180# temp102 vdd w_490_n166# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1009 vdd temp107 temp108 w_670_n220# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1010 a_348_n227# b1 vdd w_301_n233# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1011 gnd b2 a_542_n346# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1012 a_41_n338# a0 mid_s0 Gnd nfet w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1013 p1_inv b1 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1014 c2 a_546_n208# vdd w_490_n166# pfet w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1015 vdd mid_s1 a_344_n318# w_360_n325# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1016 a_248_n261# temp100 gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1017 gnd a0 a_101_n259# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1018 a_546_n208# temp102 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1019 a_789_n183# g1_inv gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1020 vdd g0_inv c1 w_162_n207# pfet w=20 l=2
+  ad=0 pd=0 as=260 ps=106
M1021 vdd a0 g0_inv w_88_n227# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1022 temp100 a_199_n249# vdd w_162_n207# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1023 vdd a_387_n246# temp102 w_375_n226# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1024 c2 a_546_n208# gnd Gnd nfet w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1025 a_135_n221# b0 vdd w_88_n227# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1026 gnd a0 p0_inv Gnd nfet w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1027 temp105 p2_inv a_786_n260# w_773_n266# pfet w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1028 gnd p2_inv temp105 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1029 a_503_n198# temp103 gnd Gnd nfet w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1030 temp100 a_199_n249# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1031 a_410_n252# c0 a_387_n246# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1032 vdd p0_inv a_461_n228# w_448_n234# pfet w=40 l=2
+  ad=0 pd=0 as=320 ps=96
M1033 gnd p0_inv temp101 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1034 vdd g1_inv temp104 w_490_n166# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1035 a_837_n246# c1 a_837_n284# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=160 ps=56
M1036 a_744_n230# g2_inv temp108 Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1037 temp108 g2_inv vdd w_670_n220# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 a_789_n193# g1_inv vdd w_783_n206# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1039 vdd temp101 a_387_n246# w_375_n226# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1040 s2 c2 a_632_n320# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1041 a_101_n259# b0 g0_inv Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1042 c1 temp100 vdd w_162_n207# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 temp103 a_398_n161# vdd w_418_n146# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1044 c0 mid_s0 s0 w_186_n314# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1045 gnd a2 a_602_n267# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1046 g0_inv b0 vdd w_88_n227# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 gnd p2_inv a_789_n183# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 mid_s2 a_542_n346# a2 Gnd nfet w=10 l=2
+  ad=70 pd=34 as=50 ps=30
M1049 gnd mid_s2 a_632_n320# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gnd a1 a_314_n265# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1051 s1 c1 a_344_n318# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1052 mid_s0 b0 a0 w_30_n314# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1053 p0_inv b0 gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 a_786_n260# p1_inv vdd w_773_n266# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 a_426_n161# g0_inv vdd w_418_n146# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1056 mid_s1 a_254_n344# a1 Gnd nfet w=10 l=2
+  ad=70 pd=34 as=50 ps=30
M1057 temp105 p1_inv gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 gnd mid_s1 a_344_n318# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 vdd mid_s0 a_131_n312# w_147_n319# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1060 a_542_n346# a2 mid_s2 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 gnd b0 a_41_n338# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 a_701_n212# temp108 a_681_n239# w_670_n220# pfet w=40 l=2
+  ad=320 pd=96 as=200 ps=90
M1063 a_461_n228# p1_inv temp101 w_448_n234# pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1064 b0 a0 mid_s0 w_30_n314# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1065 temp101 p1_inv gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 temp104 temp103 vdd w_490_n166# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_254_n344# a1 mid_s1 Gnd nfet w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1068 a_837_n284# temp105 gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 vdd a_681_n239# c3 w_670_n220# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1070 s0 c0 a_131_n312# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1071 s2 c2 mid_s2 w_687_n322# pfet w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1072 vdd b0 a_41_n338# w_70_n319# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1073 a_199_n221# p0_inv vdd w_162_n207# pfet w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1074 a_387_n246# c0 vdd w_375_n226# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 vdd c1 a_837_n246# w_824_n252# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1076 a_398_n161# g0_inv gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1077 vdd temp106 a_701_n212# w_670_n220# pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 a_789_n183# p2_inv a_789_n193# w_783_n206# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1079 temp107 a_789_n183# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1080 gnd a_681_n239# c3 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1081 temp107 a_789_n183# vdd w_783_n206# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1082 a_602_n267# b2 g2_inv Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1083 mid_s2 b2 a2 w_531_n322# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1084 a_199_n249# c0_inv a_199_n221# w_162_n207# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1085 s1 c1 mid_s1 w_399_n320# pfet w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1086 a_314_n265# b1 g1_inv Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1087 mid_s1 b1 a1 w_243_n320# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1088 vdd a2 g2_inv w_589_n235# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1089 b2 a2 mid_s2 w_531_n322# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1090 temp106 a_837_n246# vdd w_824_n252# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1091 c2 a_632_n320# s2 Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 vdd a1 g1_inv w_301_n233# pfet w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1093 vdd b2 a_542_n346# w_571_n327# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1094 b1 a1 mid_s1 w_243_n320# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1095 a_681_n239# temp108 gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1096 p2_inv a2 a_636_n229# w_589_n235# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1097 c1 a_344_n318# s1 Gnd nfet w=10 l=2
+  ad=150 pd=80 as=0 ps=0
M1098 vdd b1 a_254_n344# w_283_n325# pfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1099 gnd a2 p2_inv Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 a_398_n161# p1_inv a_426_n161# w_418_n146# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1101 temp103 a_398_n161# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1102 a_546_n208# temp104 a_546_n180# w_490_n166# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1103 a_199_n249# p0_inv gnd Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1104 temp106 a_837_n246# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1105 p1_inv a1 a_348_n227# w_301_n233# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1106 gnd a1 p1_inv Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 a_837_n246# temp105 vdd w_824_n252# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 c1 g0_inv a_248_n261# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 gnd b1 a_254_n344# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 gnd temp106 a_681_n239# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 gnd temp104 a_546_n208# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 c0_inv c0 vdd w_162_n207# pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1113 gnd mid_s0 a_131_n312# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 gnd p1_inv a_398_n161# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1115 gnd c0_inv a_199_n249# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 c0 a_131_n312# s0 Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1117 g2_inv b2 vdd w_589_n235# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 c2 mid_s2 s2 w_687_n322# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 c0_inv c0 gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1120 p0_inv a0 a_135_n221# w_88_n227# pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1121 g1_inv b1 vdd w_301_n233# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 temp104 g1_inv a_503_n198# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1123 c1 mid_s1 s1 w_399_n320# pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 p1_inv a_398_n161# 0.17fF
C1 mid_s0 a0 0.40fF
C2 a_837_n246# c1 0.10fF
C3 g1_inv temp104 0.18fF
C4 a_542_n346# a2 0.10fF
C5 b2 w_571_n327# 0.07fF
C6 c0 a1 0.01fF
C7 c0_inv a_199_n249# 0.17fF
C8 b0 mid_s0 0.25fF
C9 vdd temp107 0.84fF
C10 temp104 temp102 0.24fF
C11 w_243_n320# b1 0.10fF
C12 p1_inv a_387_n246# 0.01fF
C13 temp101 temp102 0.01fF
C14 vdd w_773_n266# 0.02fF
C15 w_399_n320# c1 0.24fF
C16 temp106 a_786_n260# 0.01fF
C17 vdd w_571_n327# 0.11fF
C18 p1_inv w_773_n266# 0.06fF
C19 w_375_n226# p0_inv 0.01fF
C20 g2_inv temp107 0.26fF
C21 w_399_n320# c0 0.01fF
C22 g0_inv p0_inv 0.05fF
C23 w_490_n166# g1_inv 0.09fF
C24 a_426_n161# g1_inv 0.03fF
C25 temp101 w_448_n234# 0.05fF
C26 g0_inv w_418_n146# 0.06fF
C27 a_41_n338# a0 0.10fF
C28 g1_inv b1 0.26fF
C29 w_670_n220# temp107 0.07fF
C30 b2 w_589_n235# 0.14fF
C31 w_490_n166# temp102 0.06fF
C32 w_301_n233# vdd 0.12fF
C33 temp106 temp105 0.01fF
C34 w_186_n314# c0 0.24fF
C35 gnd w_375_n226# 0.01fF
C36 b0 a_41_n338# 0.06fF
C37 w_70_n319# vdd 0.11fF
C38 c2 s2 0.35fF
C39 gnd g0_inv 0.09fF
C40 w_301_n233# p1_inv 0.02fF
C41 c2 w_490_n166# 0.02fF
C42 mid_s1 b1 0.25fF
C43 w_283_n325# b1 0.07fF
C44 g0_inv c1 0.10fF
C45 vdd w_589_n235# 0.12fF
C46 temp103 g1_inv 0.32fF
C47 gnd a_789_n183# 0.04fF
C48 gnd p0_inv 0.61fF
C49 w_375_n226# c0 0.07fF
C50 w_162_n207# a_199_n249# 0.09fF
C51 b2 vdd 0.19fF
C52 temp103 temp102 0.00fF
C53 p2_inv g1_inv 0.28fF
C54 g0_inv c0 0.07fF
C55 a2 w_589_n235# 0.44fF
C56 s2 w_687_n322# 0.17fF
C57 p0_inv c1 0.17fF
C58 mid_s0 w_147_n319# 0.07fF
C59 gnd mid_s2 0.22fF
C60 b2 p1_inv 0.19fF
C61 b0 w_70_n319# 0.07fF
C62 a_602_n267# b2 0.01fF
C63 vdd w_648_n327# 0.11fF
C64 g2_inv w_589_n235# 0.30fF
C65 mid_s2 c1 0.01fF
C66 b2 a2 1.02fF
C67 gnd a_546_n208# 0.04fF
C68 temp100 g0_inv 0.31fF
C69 w_186_n314# s0 0.17fF
C70 a1 b1 1.02fF
C71 c0 p0_inv 0.25fF
C72 g1_inv a_398_n161# 0.07fF
C73 g2_inv a_681_n239# 0.07fF
C74 b2 g2_inv 0.27fF
C75 w_360_n325# c0 0.02fF
C76 gnd c1 0.36fF
C77 p1_inv vdd 0.63fF
C78 a_681_n239# w_670_n220# 0.09fF
C79 temp100 p0_inv 0.00fF
C80 vdd a2 0.12fF
C81 vdd a0 0.12fF
C82 gnd c0 0.74fF
C83 mid_s2 w_531_n322# 0.18fF
C84 c2 a_632_n320# 0.10fF
C85 temp106 w_824_n252# 0.48fF
C86 p1_inv a2 0.25fF
C87 g2_inv vdd 0.07fF
C88 temp107 g1_inv 0.04fF
C89 w_162_n207# c0_inv 0.12fF
C90 c0 c1 0.12fF
C91 w_375_n226# temp101 0.07fF
C92 p2_inv temp106 0.06fF
C93 b0 vdd 0.19fF
C94 a_387_n246# temp102 0.04fF
C95 a_837_n246# w_824_n252# 0.11fF
C96 gnd a_131_n312# 0.02fF
C97 mid_s0 w_30_n314# 0.18fF
C98 w_670_n220# vdd 0.11fF
C99 g2_inv a2 0.32fF
C100 a_254_n344# w_283_n325# 0.02fF
C101 vdd w_162_n207# 0.14fF
C102 p2_inv w_783_n206# 0.07fF
C103 temp101 p0_inv 0.08fF
C104 b0 a0 0.71fF
C105 a_131_n312# c0 0.10fF
C106 g2_inv w_670_n220# 0.38fF
C107 g2_inv a_744_n230# 0.01fF
C108 a_410_n252# p1_inv 0.01fF
C109 w_301_n233# g1_inv 0.04fF
C110 a_546_n208# temp104 0.17fF
C111 gnd temp105 0.02fF
C112 a_314_n265# b1 0.01fF
C113 temp105 c1 0.25fF
C114 gnd temp101 0.02fF
C115 temp106 temp107 0.00fF
C116 a_254_n344# a1 0.10fF
C117 temp106 w_773_n266# 0.01fF
C118 p0_inv b1 0.01fF
C119 s0 c0 0.41fF
C120 mid_s0 w_186_n314# 0.10fF
C121 mid_s2 s2 0.00fF
C122 a_681_n239# g1_inv 0.00fF
C123 temp107 w_783_n206# 0.09fF
C124 c0 temp101 0.30fF
C125 w_490_n166# a_546_n208# 0.09fF
C126 gnd b1 0.05fF
C127 w_147_n319# vdd 0.11fF
C128 vdd g1_inv 0.35fF
C129 b1 c1 0.20fF
C130 temp103 w_418_n146# 0.09fF
C131 w_301_n233# a1 0.44fF
C132 p2_inv a_789_n183# 0.17fF
C133 p1_inv g1_inv 0.05fF
C134 vdd temp102 0.24fF
C135 g0_inv a_398_n161# 0.02fF
C136 vdd w_88_n227# 0.12fF
C137 vdd mid_s1 0.12fF
C138 vdd w_283_n325# 0.11fF
C139 c0 b1 0.04fF
C140 p1_inv temp102 0.06fF
C141 gnd w_824_n252# 0.01fF
C142 g2_inv g1_inv 0.00fF
C143 temp106 a_681_n239# 0.02fF
C144 vdd w_448_n234# 0.02fF
C145 a_387_n246# w_375_n226# 0.11fF
C146 w_824_n252# c1 0.07fF
C147 c2 p1_inv 0.01fF
C148 p2_inv gnd 0.14fF
C149 w_670_n220# g1_inv 0.02fF
C150 w_418_n146# a_398_n161# 0.09fF
C151 w_88_n227# a0 0.44fF
C152 a_461_n228# temp102 0.01fF
C153 b0 a_101_n259# 0.01fF
C154 p2_inv c1 0.00fF
C155 p1_inv w_448_n234# 0.47fF
C156 mid_s2 a_632_n320# 0.06fF
C157 mid_s0 gnd 0.22fF
C158 b0 w_88_n227# 0.14fF
C159 a_789_n183# temp107 0.04fF
C160 temp106 vdd 0.24fF
C161 gnd a_632_n320# 0.02fF
C162 gnd a_398_n161# 0.04fF
C163 a_387_n246# p0_inv 0.01fF
C164 vdd a1 0.12fF
C165 g0_inv a_199_n249# 0.05fF
C166 temp106 p1_inv 0.00fF
C167 w_490_n166# temp104 0.13fF
C168 p1_inv a1 0.17fF
C169 w_30_n314# a0 0.24fF
C170 mid_s0 c0 0.27fF
C171 vdd w_783_n206# 0.09fF
C172 a_199_n249# p0_inv 0.02fF
C173 gnd a_387_n246# 0.06fF
C174 temp106 g2_inv 0.02fF
C175 b0 w_30_n314# 0.10fF
C176 mid_s0 a_131_n312# 0.06fF
C177 temp106 w_670_n220# 0.06fF
C178 temp106 a_744_n230# 0.01fF
C179 a_344_n318# mid_s1 0.06fF
C180 temp105 w_824_n252# 0.07fF
C181 w_301_n233# p0_inv 0.02fF
C182 gnd a_199_n249# 0.04fF
C183 temp108 a_681_n239# 0.17fF
C184 a_387_n246# c0 0.10fF
C185 p2_inv temp105 0.17fF
C186 a_254_n344# c0 0.22fF
C187 g0_inv c0_inv 0.12fF
C188 w_243_n320# mid_s1 0.18fF
C189 p0_inv a_348_n227# 0.01fF
C190 mid_s0 s0 0.00fF
C191 vdd w_375_n226# 0.07fF
C192 c0_inv p0_inv 0.25fF
C193 g1_inv temp102 0.09fF
C194 g0_inv vdd 0.73fF
C195 temp103 w_490_n166# 0.07fF
C196 temp100 a_199_n249# 0.04fF
C197 b2 mid_s2 0.25fF
C198 p1_inv g0_inv 0.27fF
C199 c2 g1_inv 0.05fF
C200 w_243_n320# a1 0.24fF
C201 gnd a_681_n239# 0.04fF
C202 vdd p0_inv 0.09fF
C203 gnd c0_inv 0.03fF
C204 gnd b2 0.18fF
C205 temp108 g2_inv 0.36fF
C206 mid_s2 w_648_n327# 0.07fF
C207 g0_inv a0 0.38fF
C208 w_418_n146# vdd 0.09fF
C209 w_360_n325# vdd 0.11fF
C210 p1_inv p0_inv 0.42fF
C211 b2 c1 0.02fF
C212 w_773_n266# temp105 0.05fF
C213 w_448_n234# temp102 0.01fF
C214 mid_s2 vdd 0.12fF
C215 temp108 w_670_n220# 0.13fF
C216 p1_inv w_418_n146# 0.07fF
C217 b0 g0_inv 0.26fF
C218 a0 p0_inv 0.17fF
C219 gnd vdd 1.59fF
C220 temp106 g1_inv 0.00fF
C221 s1 mid_s1 0.00fF
C222 c0 c0_inv 0.04fF
C223 g1_inv a1 0.32fF
C224 mid_s2 a2 0.40fF
C225 a_461_n228# p0_inv 0.01fF
C226 vdd c1 0.12fF
C227 g0_inv w_162_n207# 0.56fF
C228 a_681_n239# c3 0.04fF
C229 gnd p1_inv 0.79fF
C230 a_602_n267# gnd 0.01fF
C231 b0 p0_inv 0.02fF
C232 gnd a2 0.14fF
C233 b2 w_531_n322# 0.10fF
C234 g1_inv w_783_n206# 0.11fF
C235 p1_inv c1 0.00fF
C236 c2 w_687_n322# 0.24fF
C237 mid_s1 a1 0.40fF
C238 a2 c1 0.04fF
C239 vdd c0 0.21fF
C240 temp103 a_398_n161# 0.04fF
C241 gnd g2_inv 0.01fF
C242 w_162_n207# p0_inv 0.06fF
C243 a_254_n344# b1 0.06fF
C244 p1_inv c0 0.06fF
C245 b0 gnd 0.05fF
C246 w_399_n320# mid_s1 0.10fF
C247 a2 w_531_n322# 0.24fF
C248 w_360_n325# a_344_n318# 0.02fF
C249 w_162_n207# c1 0.04fF
C250 g2_inv c3 0.06fF
C251 w_301_n233# b1 0.14fF
C252 a_837_n246# temp106 0.04fF
C253 s1 w_399_n320# 0.17fF
C254 w_670_n220# c3 0.02fF
C255 p2_inv w_773_n266# 0.37fF
C256 temp108 g1_inv 0.01fF
C257 gnd a_344_n318# 0.02fF
C258 w_162_n207# c0 0.07fF
C259 g0_inv g1_inv 0.05fF
C260 a_344_n318# c1 0.10fF
C261 p1_inv temp105 0.02fF
C262 w_375_n226# temp102 0.48fF
C263 temp100 w_162_n207# 0.09fF
C264 p1_inv temp101 0.33fF
C265 a_789_n183# g1_inv 0.06fF
C266 g0_inv w_88_n227# 0.30fF
C267 g1_inv p0_inv 0.06fF
C268 a_248_n261# p0_inv 0.00fF
C269 a_542_n346# w_571_n327# 0.02fF
C270 w_418_n146# g1_inv 0.01fF
C271 temp102 p0_inv 0.06fF
C272 g2_inv a_636_n229# 0.01fF
C273 vdd w_490_n166# 0.11fF
C274 w_88_n227# p0_inv 0.02fF
C275 a_546_n208# g1_inv 0.04fF
C276 vdd b1 0.19fF
C277 gnd g1_inv 0.09fF
C278 g0_inv a_199_n221# 0.01fF
C279 w_360_n325# mid_s1 0.07fF
C280 p2_inv w_589_n235# 0.02fF
C281 p1_inv b1 0.02fF
C282 a_546_n208# temp102 0.02fF
C283 temp106 temp108 0.24fF
C284 w_448_n234# p0_inv 0.07fF
C285 gnd temp102 0.11fF
C286 a_135_n221# g0_inv 0.01fF
C287 c2 mid_s2 0.27fF
C288 p2_inv b2 0.02fF
C289 gnd mid_s1 0.22fF
C290 c2 a_546_n208# 0.04fF
C291 a_701_n212# g1_inv 0.01fF
C292 temp103 vdd 0.84fF
C293 vdd w_824_n252# 0.07fF
C294 mid_s1 c1 0.27fF
C295 c2 c1 0.03fF
C296 a_131_n312# w_147_n319# 0.02fF
C297 a1 p0_inv 0.05fF
C298 c0 temp102 0.00fF
C299 p2_inv vdd 0.56fF
C300 b2 a_542_n346# 0.06fF
C301 mid_s2 w_687_n322# 0.10fF
C302 mid_s1 c0 0.05fF
C303 w_283_n325# c0 0.01fF
C304 a_789_n183# w_783_n206# 0.09fF
C305 s1 c1 0.35fF
C306 w_70_n319# a_41_n338# 0.02fF
C307 p2_inv p1_inv 0.28fF
C308 a_632_n320# w_648_n327# 0.02fF
C309 mid_s0 vdd 0.12fF
C310 p2_inv a2 0.17fF
C311 a_503_n198# g1_inv 0.01fF
C312 gnd temp106 0.11fF
C313 p2_inv g2_inv 0.03fF
C314 s1 c0 0.01fF
C315 temp106 c1 0.00fF
C316 a1 c1 0.25fF
C317 a_503_n198# temp102 0.01fF
C318 a_837_n246# gnd 0.06fF
C319 s2 Gnd 0.43fF
C320 a_632_n320# Gnd 0.38fF
C321 a_542_n346# Gnd 0.38fF
C322 c2 Gnd 0.75fF
C323 mid_s2 Gnd 1.09fF
C324 s1 Gnd 0.43fF
C325 a_344_n318# Gnd 0.38fF
C326 a_254_n344# Gnd 0.38fF
C327 mid_s1 Gnd 1.09fF
C328 s0 Gnd 0.43fF
C329 a_131_n312# Gnd 0.38fF
C330 a_41_n338# Gnd 0.38fF
C331 mid_s0 Gnd 1.09fF
C332 a_837_n246# Gnd 0.18fF
C333 temp105 Gnd 0.07fF
C334 c3 Gnd 0.04fF
C335 a_681_n239# Gnd 0.18fF
C336 p2_inv Gnd 2.82fF
C337 a2 Gnd 1.34fF
C338 b2 Gnd 1.19fF
C339 gnd Gnd 4.38fF
C340 g2_inv Gnd 1.41fF
C341 temp106 Gnd 0.14fF
C342 temp108 Gnd 0.17fF
C343 vdd Gnd 7.01fF
C344 a_789_n183# Gnd 0.18fF
C345 temp107 Gnd 0.32fF
C346 a_546_n208# Gnd 0.18fF
C347 a_387_n246# Gnd 0.18fF
C348 temp101 Gnd 0.31fF
C349 c1 Gnd 0.07fF
C350 temp100 Gnd 0.19fF
C351 a1 Gnd 0.15fF
C352 b1 Gnd 0.07fF
C353 a_199_n249# Gnd 0.18fF
C354 c0_inv Gnd 0.09fF
C355 p0_inv Gnd 1.47fF
C356 c0 Gnd 0.24fF
C357 a0 Gnd 1.78fF
C358 b0 Gnd 1.19fF
C359 g0_inv Gnd 3.26fF
C360 p1_inv Gnd 5.51fF
C361 temp104 Gnd 0.28fF
C362 temp102 Gnd 0.54fF
C363 g1_inv Gnd 1.56fF
C364 a_398_n161# Gnd 0.02fF
C365 temp103 Gnd 0.49fF
C366 w_687_n322# Gnd 1.06fF
C367 w_648_n327# Gnd 0.84fF
C368 w_571_n327# Gnd 0.84fF
C369 w_531_n322# Gnd 1.06fF
C370 w_399_n320# Gnd 1.06fF
C371 w_360_n325# Gnd 0.84fF
C372 w_283_n325# Gnd 0.84fF
C373 w_243_n320# Gnd 0.42fF
C374 w_186_n314# Gnd 1.06fF
C375 w_147_n319# Gnd 0.84fF
C376 w_70_n319# Gnd 0.84fF
C377 w_30_n314# Gnd 1.06fF
C378 w_824_n252# Gnd 1.82fF
C379 w_773_n266# Gnd 1.78fF
C380 w_783_n206# Gnd 2.40fF
C381 w_670_n220# Gnd 2.00fF
C382 w_589_n235# Gnd 1.04fF
C383 w_448_n234# Gnd 1.78fF
C384 w_375_n226# Gnd 1.43fF
C385 w_301_n233# Gnd 0.19fF
C386 w_162_n207# Gnd 1.14fF
C387 w_88_n227# Gnd 1.09fF
C388 w_490_n166# Gnd 3.75fF
C389 w_418_n146# Gnd 2.40fF