* SPICE3 file created from CLA1.ext - technology: scmos
* Adds 1 bit and generates s0 and c1
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.option scale=0.09u
.global gnd vdd

M1000 s0 mid_s0 c0 w_n91_n115# CMOSP w=20 l=2
+  ad=140 pd=54 as=100 ps=50
M1001 a_66_n170# a0 gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=600 ps=340
M1002 b0_inv a0 mid_s0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=70 ps=34
M1003 a_32_n217# a0 vdd w_n45_n202# CMOSP w=40 l=2
+  ad=320 pd=96 as=1200 ps=580
M1004 a_17_n116# c0_inv a_17_n88# w_n20_n74# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1005 mid_s0 b0_inv a0 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1006 g0_inv a0 vdd w_n45_n202# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1007 vdd g0_inv c1 w_n20_n74# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1008 a_n80_n139# c0 s0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=70 ps=34
M1009 b0_inv b0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 gnd b0 p0_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1011 a_17_n88# p0_inv vdd w_n20_n74# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 temp100 a_17_n116# vdd w_n20_n74# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1013 c0_inv c0 vdd w_n20_n74# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1014 b0_inv b0 vdd w_n45_n202# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1015 gnd c0_inv a_17_n116# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1016 c0_inv c0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1017 c1 temp100 vdd w_n20_n74# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 s0 a_n80_n139# c0 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1019 p0_inv a0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 c1 g0_inv a_66_n128# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=160 ps=56
M1021 mid_s0 c0 s0 w_n91_n115# CMOSP w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1022 a_17_n116# p0_inv gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 a_n80_n139# mid_s0 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 g0_inv b0 a_66_n170# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1025 temp100 a_17_n116# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1026 p0_inv b0 a_32_n217# w_n45_n202# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1027 a_n80_n139# mid_s0 vdd w_n91_n115# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1028 a_66_n128# temp100 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 b0 a0 mid_s0 w_n45_n202# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1030 vdd b0 g0_inv w_n45_n202# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 mid_s0 b0 a0 w_n45_n202# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
C0 b0_inv p0_inv 0.01fF
C1 a_n80_n139# gnd 0.18fF
C2 b0 p0_inv 0.30fF
C3 mid_s0 s0 0.00fF
C4 a0 p0_inv 0.05fF
C5 w_n20_n74# a_17_n116# 0.09fF
C6 c0 gnd 0.02fF
C7 w_n20_n74# vdd 0.14fF
C8 vdd mid_s0 0.23fF
C9 c0_inv p0_inv 0.25fF
C10 w_n20_n74# c1 0.04fF
C11 w_n91_n115# mid_s0 0.27fF
C12 w_n45_n202# mid_s0 0.17fF
C13 b0 mid_s0 0.00fF
C14 a0 mid_s0 0.42fF
C15 w_n20_n74# c0_inv 0.12fF
C16 g0_inv p0_inv 0.24fF
C17 c0 s0 0.34fF
C18 a_n80_n139# w_n91_n115# 0.02fF
C19 a_17_n116# temp100 0.04fF
C20 vdd c0 0.09fF
C21 a_17_n116# gnd 0.04fF
C22 w_n91_n115# c0 0.10fF
C23 w_n20_n74# g0_inv 0.07fF
C24 b0_inv gnd 0.19fF
C25 b0 gnd 0.02fF
C26 g0_inv a_66_n170# 0.01fF
C27 a0 gnd 0.02fF
C28 c0_inv c0 0.04fF
C29 w_n20_n74# p0_inv 0.06fF
C30 a0 a_32_n217# 0.01fF
C31 vdd s0 0.07fF
C32 w_n91_n115# s0 0.17fF
C33 w_n91_n115# vdd 0.02fF
C34 w_n45_n202# vdd 0.15fF
C35 g0_inv temp100 0.24fF
C36 g0_inv gnd 0.21fF
C37 b0 vdd 0.06fF
C38 w_n45_n202# b0_inv 0.02fF
C39 a0 vdd 0.00fF
C40 b0 w_n45_n202# 0.87fF
C41 a_17_n116# c0_inv 0.17fF
C42 a0 w_n45_n202# 0.37fF
C43 b0 b0_inv 0.13fF
C44 a0 b0_inv 0.09fF
C45 gnd p0_inv 0.67fF
C46 b0 a0 0.67fF
C47 a_n80_n139# mid_s0 0.23fF
C48 w_n20_n74# c0 0.09fF
C49 w_n20_n74# temp100 0.09fF
C50 c0 mid_s0 0.20fF
C51 mid_s0 gnd 0.18fF
C52 g0_inv c1 0.10fF
C53 w_n45_n202# g0_inv 0.04fF
C54 b0 g0_inv 0.11fF
C55 a_17_n116# p0_inv 0.02fF
C56 a0 g0_inv 0.00fF
C57 w_n45_n202# p0_inv 0.02fF
C58 a_n80_n139# c0 0.05fF
C59 b0 Gnd 0.15fF
C60 a0 Gnd 0.47fF
C61 b0_inv Gnd 0.23fF
C62 c1 Gnd 0.06fF
C63 g0_inv Gnd 0.17fF
C64 temp100 Gnd 0.16fF
C65 a_17_n116# Gnd 0.18fF
C66 a_n80_n139# Gnd 0.73fF
C67 s0 Gnd 5.30fF
C68 gnd Gnd 1.32fF
C69 mid_s0 Gnd 0.21fF
C70 vdd Gnd 0.03fF
C71 c0_inv Gnd 0.01fF
C72 p0_inv Gnd 0.41fF
C73 c0 Gnd 0.63fF
C74 w_n45_n202# Gnd 1.00fF
C75 w_n91_n115# Gnd 1.96fF
C76 w_n20_n74# Gnd 4.13fF

Vdd vdd gnd 'SUPPLY'
Va0 a0 gnd 0
Vb0 b0 gnd 1.8
Vc0 c0 gnd 1.8

.tran 100ps 400ns
.measure tran a0 FIND v(a0) AT=200ns
.measure tran b0 FIND v(b0) AT=200ns
.measure tran c0 FIND v(c0) AT=200ns
.measure tran s0 FIND v(s0) AT=200ns
.measure tran c1 FIND v(c1) AT=200ns

.control
set hcopypscolor = 0
set color0=white 
set color1=black 

run

set curplottitle="2023112005_1_bit_adder"

plot a0, b0+2, c0+4, s0+6, c1+8
.endc