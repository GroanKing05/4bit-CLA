magic
tech scmos
timestamp 1731430887
<< nwell >>
rect 233 -707 265 -688
rect 233 -713 287 -707
rect 235 -741 287 -713
rect 305 -723 382 -701
rect 305 -733 400 -723
rect -63 -762 -29 -742
rect -97 -794 -29 -762
rect -23 -764 35 -742
rect -23 -774 84 -764
rect 150 -768 184 -748
rect 212 -761 246 -755
rect 1 -794 84 -774
rect 29 -796 84 -794
rect 116 -800 184 -768
rect 190 -787 246 -761
rect 190 -793 215 -787
rect 263 -801 297 -749
rect 348 -753 400 -733
rect 376 -755 400 -753
rect 438 -770 472 -750
rect 503 -755 580 -733
rect 620 -739 652 -720
rect 404 -802 472 -770
rect 485 -765 580 -755
rect 598 -745 652 -739
rect 485 -785 537 -765
rect 598 -773 650 -745
rect 799 -774 833 -754
rect 485 -787 509 -785
rect 588 -833 622 -781
rect 639 -793 673 -787
rect 639 -819 695 -793
rect 765 -806 833 -774
rect 849 -757 883 -752
rect 849 -763 920 -757
rect 849 -789 942 -763
rect 976 -777 1010 -757
rect 976 -779 1044 -777
rect 849 -804 883 -789
rect 917 -795 942 -789
rect 957 -783 1044 -779
rect 957 -809 1065 -783
rect 957 -811 982 -809
rect 1041 -815 1065 -809
rect 1076 -789 1110 -767
rect 1076 -819 1129 -789
rect 670 -825 695 -819
rect 1104 -821 1129 -819
rect 1135 -821 1169 -789
rect -155 -881 -122 -849
rect -115 -886 -83 -860
rect -38 -886 -6 -860
rect 1 -881 34 -849
rect 58 -887 91 -855
rect 98 -892 130 -866
rect 175 -892 207 -866
rect 214 -887 247 -855
rect 346 -889 379 -857
rect 386 -894 418 -868
rect 463 -894 495 -868
rect 502 -889 535 -857
rect 707 -893 740 -861
rect 747 -898 779 -872
rect 824 -898 856 -872
rect 863 -893 896 -861
rect 948 -932 980 -864
rect 1057 -893 1109 -859
<< ntransistor >>
rect 217 -702 227 -700
rect 213 -720 223 -718
rect 213 -730 223 -728
rect -12 -790 -10 -780
rect -86 -826 -84 -806
rect -76 -826 -74 -806
rect -52 -816 -50 -806
rect -42 -816 -40 -806
rect 12 -816 14 -806
rect 22 -816 24 -806
rect 40 -812 42 -802
rect 61 -828 63 -808
rect 71 -828 73 -808
rect 316 -765 318 -745
rect 326 -765 328 -745
rect 658 -734 668 -732
rect 359 -775 361 -765
rect 369 -775 371 -765
rect 387 -771 389 -761
rect 202 -809 204 -799
rect 127 -832 129 -812
rect 137 -832 139 -812
rect 161 -822 163 -812
rect 171 -822 173 -812
rect 223 -819 225 -799
rect 233 -819 235 -799
rect 662 -752 672 -750
rect 662 -762 672 -760
rect 274 -823 276 -813
rect 284 -823 286 -813
rect 496 -803 498 -793
rect 557 -797 559 -777
rect 567 -797 569 -777
rect 514 -807 516 -797
rect 524 -807 526 -797
rect 415 -834 417 -814
rect 425 -834 427 -814
rect 449 -824 451 -814
rect 459 -824 461 -814
rect -77 -874 -67 -872
rect -54 -874 -44 -872
rect 136 -880 146 -878
rect 159 -880 169 -878
rect -144 -898 -142 -888
rect -135 -898 -133 -888
rect 12 -898 14 -888
rect 21 -898 23 -888
rect 599 -855 601 -845
rect 609 -855 611 -845
rect 650 -851 652 -831
rect 660 -851 662 -831
rect 681 -841 683 -831
rect 776 -838 778 -818
rect 786 -838 788 -818
rect 810 -828 812 -818
rect 820 -828 822 -818
rect 860 -826 862 -816
rect 870 -826 872 -816
rect 897 -821 899 -801
rect 907 -821 909 -801
rect 928 -811 930 -801
rect 969 -827 971 -817
rect 987 -831 989 -821
rect 997 -831 999 -821
rect 1021 -841 1023 -821
rect 1031 -841 1033 -821
rect 1052 -831 1054 -821
rect 1087 -841 1089 -831
rect 1097 -841 1099 -831
rect 1115 -837 1117 -827
rect 1146 -853 1148 -833
rect 1156 -853 1158 -833
rect 424 -882 434 -880
rect 447 -882 457 -880
rect 69 -904 71 -894
rect 78 -904 80 -894
rect 225 -904 227 -894
rect 234 -904 236 -894
rect 785 -886 795 -884
rect 808 -886 818 -884
rect 357 -906 359 -896
rect 366 -906 368 -896
rect 513 -906 515 -896
rect 522 -906 524 -896
rect 1121 -872 1131 -870
rect 992 -877 1012 -875
rect 1121 -882 1131 -880
rect 992 -887 1012 -885
rect 718 -910 720 -900
rect 727 -910 729 -900
rect 874 -910 876 -900
rect 883 -910 885 -900
rect 992 -911 1012 -909
rect 992 -921 1012 -919
<< ptransistor >>
rect 239 -702 259 -700
rect 241 -720 281 -718
rect 316 -727 318 -707
rect 326 -727 328 -707
rect 241 -730 281 -728
rect -86 -788 -84 -768
rect -76 -788 -74 -768
rect -52 -788 -50 -748
rect -42 -788 -40 -748
rect -12 -768 -10 -748
rect 12 -788 14 -748
rect 22 -788 24 -748
rect 40 -790 42 -770
rect 61 -790 63 -770
rect 71 -790 73 -770
rect 127 -794 129 -774
rect 137 -794 139 -774
rect 161 -794 163 -754
rect 171 -794 173 -754
rect 202 -787 204 -767
rect 223 -781 225 -761
rect 233 -781 235 -761
rect 274 -795 276 -755
rect 284 -795 286 -755
rect 359 -747 361 -707
rect 369 -747 371 -707
rect 387 -749 389 -729
rect 626 -734 646 -732
rect 415 -796 417 -776
rect 425 -796 427 -776
rect 449 -796 451 -756
rect 459 -796 461 -756
rect 496 -781 498 -761
rect 514 -779 516 -739
rect 524 -779 526 -739
rect 557 -759 559 -739
rect 567 -759 569 -739
rect 604 -752 644 -750
rect 604 -762 644 -760
rect 599 -827 601 -787
rect 609 -827 611 -787
rect 650 -813 652 -793
rect 660 -813 662 -793
rect 681 -819 683 -799
rect 776 -800 778 -780
rect 786 -800 788 -780
rect 810 -800 812 -760
rect 820 -800 822 -760
rect 860 -798 862 -758
rect 870 -798 872 -758
rect 897 -783 899 -763
rect 907 -783 909 -763
rect 928 -789 930 -769
rect -144 -875 -142 -855
rect -135 -875 -133 -855
rect -109 -874 -89 -872
rect -32 -874 -12 -872
rect 12 -875 14 -855
rect 21 -875 23 -855
rect 69 -881 71 -861
rect 78 -881 80 -861
rect 104 -880 124 -878
rect 181 -880 201 -878
rect 225 -881 227 -861
rect 234 -881 236 -861
rect 969 -805 971 -785
rect 987 -803 989 -763
rect 997 -803 999 -763
rect 1021 -803 1023 -783
rect 1031 -803 1033 -783
rect 1052 -809 1054 -789
rect 1087 -813 1089 -773
rect 1097 -813 1099 -773
rect 1115 -815 1117 -795
rect 1146 -815 1148 -795
rect 1156 -815 1158 -795
rect 357 -883 359 -863
rect 366 -883 368 -863
rect 392 -882 412 -880
rect 469 -882 489 -880
rect 513 -883 515 -863
rect 522 -883 524 -863
rect 718 -887 720 -867
rect 727 -887 729 -867
rect 753 -886 773 -884
rect 830 -886 850 -884
rect 874 -887 876 -867
rect 883 -887 885 -867
rect 1063 -872 1103 -870
rect 954 -877 974 -875
rect 1063 -882 1103 -880
rect 954 -887 974 -885
rect 954 -911 974 -909
rect 954 -921 974 -919
<< ndiffusion >>
rect 217 -699 223 -695
rect 217 -700 227 -699
rect 217 -703 227 -702
rect 221 -707 227 -703
rect 217 -717 223 -713
rect 213 -718 223 -717
rect 213 -722 223 -720
rect 213 -726 219 -722
rect 213 -728 223 -726
rect 213 -731 223 -730
rect 217 -735 223 -731
rect -17 -786 -12 -780
rect -13 -790 -12 -786
rect -10 -784 -9 -780
rect -10 -790 -5 -784
rect -87 -810 -86 -806
rect -91 -826 -86 -810
rect -84 -826 -76 -806
rect -74 -822 -69 -806
rect -57 -812 -52 -806
rect -53 -816 -52 -812
rect -50 -810 -48 -806
rect -44 -810 -42 -806
rect -50 -816 -42 -810
rect -40 -812 -35 -806
rect -40 -816 -39 -812
rect 7 -812 12 -806
rect 11 -816 12 -812
rect 14 -810 16 -806
rect 20 -810 22 -806
rect 14 -816 22 -810
rect 24 -812 29 -806
rect 35 -808 40 -802
rect 39 -812 40 -808
rect 42 -806 43 -802
rect 42 -812 47 -806
rect 24 -816 25 -812
rect -74 -826 -73 -822
rect 56 -824 61 -808
rect 60 -828 61 -824
rect 63 -828 71 -808
rect 73 -812 74 -808
rect 311 -761 316 -745
rect 315 -765 316 -761
rect 318 -765 326 -745
rect 328 -749 329 -745
rect 328 -765 333 -749
rect 662 -731 668 -727
rect 658 -732 668 -731
rect 658 -735 668 -734
rect 658 -739 664 -735
rect 354 -771 359 -765
rect 358 -775 359 -771
rect 361 -769 363 -765
rect 367 -769 369 -765
rect 361 -775 369 -769
rect 371 -771 376 -765
rect 382 -767 387 -761
rect 386 -771 387 -767
rect 389 -765 390 -761
rect 389 -771 394 -765
rect 371 -775 372 -771
rect 201 -803 202 -799
rect 197 -809 202 -803
rect 204 -805 209 -799
rect 204 -809 205 -805
rect 222 -803 223 -799
rect 73 -828 78 -812
rect 126 -816 127 -812
rect 122 -832 127 -816
rect 129 -832 137 -812
rect 139 -828 144 -812
rect 156 -818 161 -812
rect 160 -822 161 -818
rect 163 -816 165 -812
rect 169 -816 171 -812
rect 163 -822 171 -816
rect 173 -818 178 -812
rect 173 -822 174 -818
rect 218 -819 223 -803
rect 225 -819 233 -799
rect 235 -815 240 -799
rect 662 -749 668 -745
rect 662 -750 672 -749
rect 662 -754 672 -752
rect 666 -758 672 -754
rect 662 -760 672 -758
rect 662 -763 672 -762
rect 662 -767 668 -763
rect 235 -819 236 -815
rect 269 -819 274 -813
rect 273 -823 274 -819
rect 276 -817 278 -813
rect 282 -817 284 -813
rect 276 -823 284 -817
rect 286 -819 291 -813
rect 495 -797 496 -793
rect 491 -803 496 -797
rect 498 -799 503 -793
rect 556 -781 557 -777
rect 552 -797 557 -781
rect 559 -797 567 -777
rect 569 -793 574 -777
rect 569 -797 570 -793
rect 498 -803 499 -799
rect 509 -803 514 -797
rect 513 -807 514 -803
rect 516 -801 518 -797
rect 522 -801 524 -797
rect 516 -807 524 -801
rect 526 -803 531 -797
rect 526 -807 527 -803
rect 286 -823 287 -819
rect 414 -818 415 -814
rect 139 -832 140 -828
rect 410 -834 415 -818
rect 417 -834 425 -814
rect 427 -830 432 -814
rect 444 -820 449 -814
rect 448 -824 449 -820
rect 451 -818 453 -814
rect 457 -818 459 -814
rect 451 -824 459 -818
rect 461 -820 466 -814
rect 461 -824 462 -820
rect 427 -834 428 -830
rect 775 -822 776 -818
rect -77 -871 -71 -867
rect -77 -872 -67 -871
rect -47 -871 -44 -867
rect -54 -872 -44 -871
rect -77 -875 -67 -874
rect -73 -879 -67 -875
rect -54 -875 -44 -874
rect -54 -879 -48 -875
rect 594 -851 599 -845
rect 136 -877 142 -873
rect 136 -878 146 -877
rect 166 -877 169 -873
rect 159 -878 169 -877
rect -145 -892 -144 -888
rect -149 -898 -144 -892
rect -142 -892 -140 -888
rect -136 -892 -135 -888
rect -142 -898 -135 -892
rect -133 -894 -128 -888
rect -133 -898 -132 -894
rect 7 -894 12 -888
rect 11 -898 12 -894
rect 14 -892 15 -888
rect 19 -892 21 -888
rect 14 -898 21 -892
rect 23 -892 24 -888
rect 23 -898 28 -892
rect 136 -881 146 -880
rect 140 -885 146 -881
rect 159 -881 169 -880
rect 159 -885 165 -881
rect 598 -855 599 -851
rect 601 -849 603 -845
rect 607 -849 609 -845
rect 601 -855 609 -849
rect 611 -851 616 -845
rect 645 -847 650 -831
rect 649 -851 650 -847
rect 652 -851 660 -831
rect 662 -835 663 -831
rect 662 -851 667 -835
rect 676 -837 681 -831
rect 680 -841 681 -837
rect 683 -835 684 -831
rect 683 -841 688 -835
rect 771 -838 776 -822
rect 778 -838 786 -818
rect 788 -834 793 -818
rect 805 -824 810 -818
rect 809 -828 810 -824
rect 812 -822 814 -818
rect 818 -822 820 -818
rect 812 -828 820 -822
rect 822 -824 827 -818
rect 822 -828 823 -824
rect 855 -822 860 -816
rect 859 -826 860 -822
rect 862 -820 864 -816
rect 868 -820 870 -816
rect 862 -826 870 -820
rect 872 -822 877 -816
rect 892 -817 897 -801
rect 896 -821 897 -817
rect 899 -821 907 -801
rect 909 -805 910 -801
rect 909 -821 914 -805
rect 923 -807 928 -801
rect 927 -811 928 -807
rect 930 -805 931 -801
rect 930 -811 935 -805
rect 968 -821 969 -817
rect 872 -826 873 -822
rect 964 -827 969 -821
rect 971 -823 976 -817
rect 971 -827 972 -823
rect 982 -827 987 -821
rect 986 -831 987 -827
rect 989 -825 991 -821
rect 995 -825 997 -821
rect 989 -831 997 -825
rect 999 -827 1004 -821
rect 999 -831 1000 -827
rect 788 -838 789 -834
rect 1016 -837 1021 -821
rect 1020 -841 1021 -837
rect 1023 -841 1031 -821
rect 1033 -825 1034 -821
rect 1033 -841 1038 -825
rect 1047 -827 1052 -821
rect 1051 -831 1052 -827
rect 1054 -825 1055 -821
rect 1054 -831 1059 -825
rect 1082 -837 1087 -831
rect 1086 -841 1087 -837
rect 1089 -835 1091 -831
rect 1095 -835 1097 -831
rect 1089 -841 1097 -835
rect 1099 -837 1104 -831
rect 1110 -833 1115 -827
rect 1114 -837 1115 -833
rect 1117 -831 1118 -827
rect 1117 -837 1122 -831
rect 1099 -841 1100 -837
rect 1141 -849 1146 -833
rect 611 -855 612 -851
rect 1145 -853 1146 -849
rect 1148 -853 1156 -833
rect 1158 -837 1159 -833
rect 1158 -853 1163 -837
rect 424 -879 430 -875
rect 424 -880 434 -879
rect 454 -879 457 -875
rect 447 -880 457 -879
rect 68 -898 69 -894
rect 64 -904 69 -898
rect 71 -898 73 -894
rect 77 -898 78 -894
rect 71 -904 78 -898
rect 80 -900 85 -894
rect 80 -904 81 -900
rect 220 -900 225 -894
rect 224 -904 225 -900
rect 227 -898 228 -894
rect 232 -898 234 -894
rect 227 -904 234 -898
rect 236 -898 237 -894
rect 424 -883 434 -882
rect 428 -887 434 -883
rect 447 -883 457 -882
rect 447 -887 453 -883
rect 785 -883 791 -879
rect 785 -884 795 -883
rect 815 -883 818 -879
rect 808 -884 818 -883
rect 236 -904 241 -898
rect 356 -900 357 -896
rect 352 -906 357 -900
rect 359 -900 361 -896
rect 365 -900 366 -896
rect 359 -906 366 -900
rect 368 -902 373 -896
rect 368 -906 369 -902
rect 508 -902 513 -896
rect 512 -906 513 -902
rect 515 -900 516 -896
rect 520 -900 522 -896
rect 515 -906 522 -900
rect 524 -900 525 -896
rect 785 -887 795 -886
rect 789 -891 795 -887
rect 808 -887 818 -886
rect 808 -891 814 -887
rect 1121 -869 1127 -865
rect 1121 -870 1131 -869
rect 992 -874 1008 -870
rect 992 -875 1012 -874
rect 992 -885 1012 -877
rect 1121 -874 1131 -872
rect 1125 -878 1131 -874
rect 1121 -880 1131 -878
rect 1121 -883 1131 -882
rect 1121 -887 1127 -883
rect 992 -888 1012 -887
rect 996 -892 1012 -888
rect 524 -906 529 -900
rect 717 -904 718 -900
rect 713 -910 718 -904
rect 720 -904 722 -900
rect 726 -904 727 -900
rect 720 -910 727 -904
rect 729 -906 734 -900
rect 729 -910 730 -906
rect 869 -906 874 -900
rect 873 -910 874 -906
rect 876 -904 877 -900
rect 881 -904 883 -900
rect 876 -910 883 -904
rect 885 -904 886 -900
rect 885 -910 890 -904
rect 992 -908 1008 -904
rect 992 -909 1012 -908
rect 992 -919 1012 -911
rect 992 -922 1012 -921
rect 996 -926 1012 -922
<< pdiffusion >>
rect 243 -699 259 -695
rect 239 -700 259 -699
rect 239 -703 259 -702
rect 239 -707 255 -703
rect 315 -711 316 -707
rect 245 -717 281 -713
rect 241 -718 281 -717
rect 241 -728 281 -720
rect 311 -727 316 -711
rect 318 -723 326 -707
rect 318 -727 320 -723
rect 324 -727 326 -723
rect 328 -711 329 -707
rect 328 -727 333 -711
rect 358 -711 359 -707
rect 241 -731 281 -730
rect 241 -735 277 -731
rect -53 -752 -52 -748
rect -87 -772 -86 -768
rect -91 -788 -86 -772
rect -84 -784 -76 -768
rect -84 -788 -82 -784
rect -78 -788 -76 -784
rect -74 -772 -73 -768
rect -74 -788 -69 -772
rect -57 -788 -52 -752
rect -50 -788 -42 -748
rect -40 -784 -35 -748
rect -13 -752 -12 -748
rect -17 -768 -12 -752
rect -10 -764 -5 -748
rect -10 -768 -9 -764
rect 11 -752 12 -748
rect -40 -788 -39 -784
rect 7 -788 12 -752
rect 14 -788 22 -748
rect 24 -784 29 -748
rect 160 -758 161 -754
rect 24 -788 25 -784
rect 39 -774 40 -770
rect 35 -790 40 -774
rect 42 -786 47 -770
rect 42 -790 43 -786
rect 60 -774 61 -770
rect 56 -790 61 -774
rect 63 -786 71 -770
rect 63 -790 65 -786
rect 69 -790 71 -786
rect 73 -774 74 -770
rect 73 -790 78 -774
rect 126 -778 127 -774
rect 122 -794 127 -778
rect 129 -790 137 -774
rect 129 -794 131 -790
rect 135 -794 137 -790
rect 139 -778 140 -774
rect 139 -794 144 -778
rect 156 -794 161 -758
rect 163 -794 171 -754
rect 173 -790 178 -754
rect 222 -765 223 -761
rect 197 -783 202 -767
rect 201 -787 202 -783
rect 204 -771 205 -767
rect 204 -787 209 -771
rect 218 -781 223 -765
rect 225 -777 233 -761
rect 225 -781 227 -777
rect 231 -781 233 -777
rect 235 -765 236 -761
rect 235 -781 240 -765
rect 173 -794 174 -790
rect 269 -791 274 -755
rect 273 -795 274 -791
rect 276 -795 284 -755
rect 286 -759 287 -755
rect 286 -795 291 -759
rect 354 -747 359 -711
rect 361 -747 369 -707
rect 371 -743 376 -707
rect 371 -747 372 -743
rect 386 -733 387 -729
rect 382 -749 387 -733
rect 389 -745 394 -729
rect 626 -731 642 -727
rect 626 -732 646 -731
rect 626 -735 646 -734
rect 630 -739 646 -735
rect 389 -749 390 -745
rect 448 -760 449 -756
rect 414 -780 415 -776
rect 410 -796 415 -780
rect 417 -792 425 -776
rect 417 -796 419 -792
rect 423 -796 425 -792
rect 427 -780 428 -776
rect 427 -796 432 -780
rect 444 -796 449 -760
rect 451 -796 459 -756
rect 461 -792 466 -756
rect 491 -777 496 -761
rect 495 -781 496 -777
rect 498 -765 499 -761
rect 498 -781 503 -765
rect 509 -775 514 -739
rect 513 -779 514 -775
rect 516 -779 524 -739
rect 526 -743 527 -739
rect 526 -779 531 -743
rect 556 -743 557 -739
rect 552 -759 557 -743
rect 559 -755 567 -739
rect 559 -759 561 -755
rect 565 -759 567 -755
rect 569 -743 570 -739
rect 569 -759 574 -743
rect 604 -749 640 -745
rect 604 -750 644 -749
rect 604 -760 644 -752
rect 604 -763 644 -762
rect 608 -767 644 -763
rect 809 -764 810 -760
rect 461 -796 462 -792
rect 775 -784 776 -780
rect 598 -791 599 -787
rect 594 -827 599 -791
rect 601 -827 609 -787
rect 611 -823 616 -787
rect 649 -797 650 -793
rect 645 -813 650 -797
rect 652 -809 660 -793
rect 652 -813 654 -809
rect 658 -813 660 -809
rect 662 -797 663 -793
rect 662 -813 667 -797
rect 680 -803 681 -799
rect 611 -827 612 -823
rect 676 -819 681 -803
rect 683 -815 688 -799
rect 771 -800 776 -784
rect 778 -796 786 -780
rect 778 -800 780 -796
rect 784 -800 786 -796
rect 788 -784 789 -780
rect 788 -800 793 -784
rect 805 -800 810 -764
rect 812 -800 820 -760
rect 822 -796 827 -760
rect 822 -800 823 -796
rect 859 -762 860 -758
rect 855 -798 860 -762
rect 862 -798 870 -758
rect 872 -794 877 -758
rect 896 -767 897 -763
rect 892 -783 897 -767
rect 899 -779 907 -763
rect 899 -783 901 -779
rect 905 -783 907 -779
rect 909 -767 910 -763
rect 909 -783 914 -767
rect 927 -773 928 -769
rect 872 -798 873 -794
rect 683 -819 684 -815
rect 923 -789 928 -773
rect 930 -785 935 -769
rect 930 -789 931 -785
rect 964 -801 969 -785
rect -149 -871 -144 -855
rect -145 -875 -144 -871
rect -142 -869 -135 -855
rect -142 -873 -140 -869
rect -136 -873 -135 -869
rect -142 -875 -135 -873
rect -133 -859 -132 -855
rect -133 -875 -128 -859
rect 11 -859 12 -855
rect -104 -871 -89 -866
rect -109 -872 -89 -871
rect -32 -871 -17 -866
rect -32 -872 -12 -871
rect -109 -875 -89 -874
rect -109 -879 -93 -875
rect -32 -875 -12 -874
rect 7 -875 12 -859
rect 14 -869 21 -855
rect 14 -873 15 -869
rect 19 -873 21 -869
rect 14 -875 21 -873
rect 23 -871 28 -855
rect 23 -875 24 -871
rect -28 -879 -12 -875
rect 64 -877 69 -861
rect 68 -881 69 -877
rect 71 -875 78 -861
rect 71 -879 73 -875
rect 77 -879 78 -875
rect 71 -881 78 -879
rect 80 -865 81 -861
rect 80 -881 85 -865
rect 224 -865 225 -861
rect 109 -877 124 -872
rect 104 -878 124 -877
rect 181 -877 196 -872
rect 181 -878 201 -877
rect 104 -881 124 -880
rect 104 -885 120 -881
rect 181 -881 201 -880
rect 220 -881 225 -865
rect 227 -875 234 -861
rect 227 -879 228 -875
rect 232 -879 234 -875
rect 227 -881 234 -879
rect 236 -877 241 -861
rect 968 -805 969 -801
rect 971 -789 972 -785
rect 971 -805 976 -789
rect 982 -799 987 -763
rect 986 -803 987 -799
rect 989 -803 997 -763
rect 999 -767 1000 -763
rect 999 -803 1004 -767
rect 1086 -777 1087 -773
rect 1020 -787 1021 -783
rect 1016 -803 1021 -787
rect 1023 -799 1031 -783
rect 1023 -803 1025 -799
rect 1029 -803 1031 -799
rect 1033 -787 1034 -783
rect 1033 -803 1038 -787
rect 1051 -793 1052 -789
rect 1047 -809 1052 -793
rect 1054 -805 1059 -789
rect 1054 -809 1055 -805
rect 1082 -813 1087 -777
rect 1089 -813 1097 -773
rect 1099 -809 1104 -773
rect 1099 -813 1100 -809
rect 1114 -799 1115 -795
rect 1110 -815 1115 -799
rect 1117 -811 1122 -795
rect 1117 -815 1118 -811
rect 1145 -799 1146 -795
rect 1141 -815 1146 -799
rect 1148 -811 1156 -795
rect 1148 -815 1150 -811
rect 1154 -815 1156 -811
rect 1158 -799 1159 -795
rect 1158 -815 1163 -799
rect 236 -881 237 -877
rect 352 -879 357 -863
rect 185 -885 201 -881
rect 356 -883 357 -879
rect 359 -877 366 -863
rect 359 -881 361 -877
rect 365 -881 366 -877
rect 359 -883 366 -881
rect 368 -867 369 -863
rect 368 -883 373 -867
rect 512 -867 513 -863
rect 397 -879 412 -874
rect 392 -880 412 -879
rect 469 -879 484 -874
rect 469 -880 489 -879
rect 392 -883 412 -882
rect 392 -887 408 -883
rect 469 -883 489 -882
rect 508 -883 513 -867
rect 515 -877 522 -863
rect 515 -881 516 -877
rect 520 -881 522 -877
rect 515 -883 522 -881
rect 524 -879 529 -863
rect 524 -883 525 -879
rect 713 -883 718 -867
rect 473 -887 489 -883
rect 717 -887 718 -883
rect 720 -881 727 -867
rect 720 -885 722 -881
rect 726 -885 727 -881
rect 720 -887 727 -885
rect 729 -871 730 -867
rect 729 -887 734 -871
rect 873 -871 874 -867
rect 758 -883 773 -878
rect 753 -884 773 -883
rect 830 -883 845 -878
rect 830 -884 850 -883
rect 753 -887 773 -886
rect 753 -891 769 -887
rect 830 -887 850 -886
rect 869 -887 874 -871
rect 876 -881 883 -867
rect 876 -885 877 -881
rect 881 -885 883 -881
rect 876 -887 883 -885
rect 885 -883 890 -867
rect 1067 -869 1103 -865
rect 1063 -870 1103 -869
rect 958 -874 974 -870
rect 954 -875 974 -874
rect 885 -887 886 -883
rect 954 -879 974 -877
rect 954 -883 970 -879
rect 954 -885 974 -883
rect 1063 -880 1103 -872
rect 1063 -883 1103 -882
rect 1063 -887 1099 -883
rect 834 -891 850 -887
rect 954 -888 974 -887
rect 958 -892 974 -888
rect 958 -908 974 -904
rect 954 -909 974 -908
rect 954 -913 974 -911
rect 954 -917 970 -913
rect 954 -919 974 -917
rect 954 -922 974 -921
rect 958 -926 974 -922
<< ndcontact >>
rect 223 -699 227 -695
rect 217 -707 221 -703
rect 213 -717 217 -713
rect 219 -726 223 -722
rect 213 -735 217 -731
rect -17 -790 -13 -786
rect -9 -784 -5 -780
rect -91 -810 -87 -806
rect -57 -816 -53 -812
rect -48 -810 -44 -806
rect -39 -816 -35 -812
rect 7 -816 11 -812
rect 16 -810 20 -806
rect 35 -812 39 -808
rect 43 -806 47 -802
rect 25 -816 29 -812
rect -73 -826 -69 -822
rect 56 -828 60 -824
rect 74 -812 78 -808
rect 311 -765 315 -761
rect 329 -749 333 -745
rect 658 -731 662 -727
rect 664 -739 668 -735
rect 354 -775 358 -771
rect 363 -769 367 -765
rect 382 -771 386 -767
rect 390 -765 394 -761
rect 372 -775 376 -771
rect 197 -803 201 -799
rect 205 -809 209 -805
rect 218 -803 222 -799
rect 122 -816 126 -812
rect 156 -822 160 -818
rect 165 -816 169 -812
rect 174 -822 178 -818
rect 668 -749 672 -745
rect 662 -758 666 -754
rect 668 -767 672 -763
rect 236 -819 240 -815
rect 269 -823 273 -819
rect 278 -817 282 -813
rect 491 -797 495 -793
rect 552 -781 556 -777
rect 570 -797 574 -793
rect 499 -803 503 -799
rect 509 -807 513 -803
rect 518 -801 522 -797
rect 527 -807 531 -803
rect 287 -823 291 -819
rect 410 -818 414 -814
rect 140 -832 144 -828
rect 444 -824 448 -820
rect 453 -818 457 -814
rect 462 -824 466 -820
rect 428 -834 432 -830
rect 771 -822 775 -818
rect -71 -871 -67 -867
rect -54 -871 -47 -867
rect -77 -879 -73 -875
rect -48 -879 -44 -875
rect 142 -877 146 -873
rect 159 -877 166 -873
rect -149 -892 -145 -888
rect -140 -892 -136 -888
rect -132 -898 -128 -894
rect 7 -898 11 -894
rect 15 -892 19 -888
rect 24 -892 28 -888
rect 136 -885 140 -881
rect 165 -885 169 -881
rect 594 -855 598 -851
rect 603 -849 607 -845
rect 645 -851 649 -847
rect 663 -835 667 -831
rect 676 -841 680 -837
rect 684 -835 688 -831
rect 805 -828 809 -824
rect 814 -822 818 -818
rect 823 -828 827 -824
rect 855 -826 859 -822
rect 864 -820 868 -816
rect 892 -821 896 -817
rect 910 -805 914 -801
rect 923 -811 927 -807
rect 931 -805 935 -801
rect 964 -821 968 -817
rect 873 -826 877 -822
rect 972 -827 976 -823
rect 982 -831 986 -827
rect 991 -825 995 -821
rect 1000 -831 1004 -827
rect 789 -838 793 -834
rect 1016 -841 1020 -837
rect 1034 -825 1038 -821
rect 1047 -831 1051 -827
rect 1055 -825 1059 -821
rect 1082 -841 1086 -837
rect 1091 -835 1095 -831
rect 1110 -837 1114 -833
rect 1118 -831 1122 -827
rect 1100 -841 1104 -837
rect 612 -855 616 -851
rect 1141 -853 1145 -849
rect 1159 -837 1163 -833
rect 430 -879 434 -875
rect 447 -879 454 -875
rect 64 -898 68 -894
rect 73 -898 77 -894
rect 81 -904 85 -900
rect 220 -904 224 -900
rect 228 -898 232 -894
rect 237 -898 241 -894
rect 424 -887 428 -883
rect 453 -887 457 -883
rect 791 -883 795 -879
rect 808 -883 815 -879
rect 352 -900 356 -896
rect 361 -900 365 -896
rect 369 -906 373 -902
rect 508 -906 512 -902
rect 516 -900 520 -896
rect 525 -900 529 -896
rect 785 -891 789 -887
rect 814 -891 818 -887
rect 1127 -869 1131 -865
rect 1008 -874 1012 -870
rect 1121 -878 1125 -874
rect 1127 -887 1131 -883
rect 992 -892 996 -888
rect 713 -904 717 -900
rect 722 -904 726 -900
rect 730 -910 734 -906
rect 869 -910 873 -906
rect 877 -904 881 -900
rect 886 -904 890 -900
rect 1008 -908 1012 -904
rect 992 -926 996 -922
<< pdcontact >>
rect 239 -699 243 -695
rect 255 -707 259 -703
rect 311 -711 315 -707
rect 241 -717 245 -713
rect 320 -727 324 -723
rect 329 -711 333 -707
rect 354 -711 358 -707
rect 277 -735 281 -731
rect -57 -752 -53 -748
rect -91 -772 -87 -768
rect -82 -788 -78 -784
rect -73 -772 -69 -768
rect -17 -752 -13 -748
rect -9 -768 -5 -764
rect 7 -752 11 -748
rect -39 -788 -35 -784
rect 156 -758 160 -754
rect 25 -788 29 -784
rect 35 -774 39 -770
rect 43 -790 47 -786
rect 56 -774 60 -770
rect 65 -790 69 -786
rect 74 -774 78 -770
rect 122 -778 126 -774
rect 131 -794 135 -790
rect 140 -778 144 -774
rect 218 -765 222 -761
rect 197 -787 201 -783
rect 205 -771 209 -767
rect 227 -781 231 -777
rect 236 -765 240 -761
rect 174 -794 178 -790
rect 269 -795 273 -791
rect 287 -759 291 -755
rect 372 -747 376 -743
rect 382 -733 386 -729
rect 642 -731 646 -727
rect 626 -739 630 -735
rect 390 -749 394 -745
rect 444 -760 448 -756
rect 410 -780 414 -776
rect 419 -796 423 -792
rect 428 -780 432 -776
rect 491 -781 495 -777
rect 499 -765 503 -761
rect 509 -779 513 -775
rect 527 -743 531 -739
rect 552 -743 556 -739
rect 561 -759 565 -755
rect 570 -743 574 -739
rect 640 -749 644 -745
rect 604 -767 608 -763
rect 805 -764 809 -760
rect 462 -796 466 -792
rect 771 -784 775 -780
rect 594 -791 598 -787
rect 645 -797 649 -793
rect 654 -813 658 -809
rect 663 -797 667 -793
rect 676 -803 680 -799
rect 612 -827 616 -823
rect 780 -800 784 -796
rect 789 -784 793 -780
rect 823 -800 827 -796
rect 855 -762 859 -758
rect 892 -767 896 -763
rect 901 -783 905 -779
rect 910 -767 914 -763
rect 923 -773 927 -769
rect 873 -798 877 -794
rect 684 -819 688 -815
rect 931 -789 935 -785
rect -149 -875 -145 -871
rect -140 -873 -136 -869
rect -132 -859 -128 -855
rect 7 -859 11 -855
rect -93 -879 -89 -875
rect 15 -873 19 -869
rect 24 -875 28 -871
rect -32 -879 -28 -875
rect 64 -881 68 -877
rect 73 -879 77 -875
rect 81 -865 85 -861
rect 220 -865 224 -861
rect 120 -885 124 -881
rect 228 -879 232 -875
rect 964 -805 968 -801
rect 972 -789 976 -785
rect 982 -803 986 -799
rect 1000 -767 1004 -763
rect 1082 -777 1086 -773
rect 1016 -787 1020 -783
rect 1025 -803 1029 -799
rect 1034 -787 1038 -783
rect 1047 -793 1051 -789
rect 1055 -809 1059 -805
rect 1100 -813 1104 -809
rect 1110 -799 1114 -795
rect 1118 -815 1122 -811
rect 1141 -799 1145 -795
rect 1150 -815 1154 -811
rect 1159 -799 1163 -795
rect 237 -881 241 -877
rect 181 -885 185 -881
rect 352 -883 356 -879
rect 361 -881 365 -877
rect 369 -867 373 -863
rect 508 -867 512 -863
rect 408 -887 412 -883
rect 516 -881 520 -877
rect 525 -883 529 -879
rect 469 -887 473 -883
rect 713 -887 717 -883
rect 722 -885 726 -881
rect 730 -871 734 -867
rect 869 -871 873 -867
rect 769 -891 773 -887
rect 877 -885 881 -881
rect 1063 -869 1067 -865
rect 954 -874 958 -870
rect 886 -887 890 -883
rect 970 -883 974 -879
rect 1099 -887 1103 -883
rect 830 -891 834 -887
rect 954 -892 958 -888
rect 954 -908 958 -904
rect 970 -917 974 -913
rect 954 -926 958 -922
<< polysilicon >>
rect 214 -702 217 -700
rect 227 -702 239 -700
rect 259 -702 262 -700
rect 316 -707 318 -703
rect 326 -707 328 -703
rect 359 -707 361 -704
rect 369 -707 371 -704
rect 210 -720 213 -718
rect 223 -720 241 -718
rect 281 -720 284 -718
rect 210 -730 213 -728
rect 223 -730 241 -728
rect 281 -730 284 -728
rect -52 -748 -50 -745
rect -42 -748 -40 -745
rect -12 -748 -10 -744
rect 316 -745 318 -727
rect 326 -745 328 -727
rect 12 -748 14 -745
rect 22 -748 24 -745
rect -86 -768 -84 -764
rect -76 -768 -74 -764
rect -12 -780 -10 -768
rect -86 -806 -84 -788
rect -76 -806 -74 -788
rect -52 -806 -50 -788
rect -42 -806 -40 -788
rect 161 -754 163 -751
rect 171 -754 173 -751
rect 40 -770 42 -767
rect 61 -770 63 -766
rect 71 -770 73 -766
rect -12 -794 -10 -790
rect 12 -806 14 -788
rect 22 -806 24 -788
rect 127 -774 129 -770
rect 137 -774 139 -770
rect 40 -802 42 -790
rect 61 -808 63 -790
rect 71 -808 73 -790
rect 274 -755 276 -752
rect 284 -755 286 -752
rect 223 -761 225 -757
rect 233 -761 235 -757
rect 202 -767 204 -763
rect 40 -815 42 -812
rect -52 -819 -50 -816
rect -42 -819 -40 -816
rect 12 -819 14 -816
rect 22 -819 24 -816
rect -86 -830 -84 -826
rect -76 -830 -74 -826
rect 127 -812 129 -794
rect 137 -812 139 -794
rect 161 -812 163 -794
rect 171 -812 173 -794
rect 202 -799 204 -787
rect 223 -799 225 -781
rect 233 -799 235 -781
rect 387 -729 389 -726
rect 359 -765 361 -747
rect 369 -765 371 -747
rect 623 -734 626 -732
rect 646 -734 658 -732
rect 668 -734 671 -732
rect 514 -739 516 -736
rect 524 -739 526 -736
rect 557 -739 559 -735
rect 567 -739 569 -735
rect 387 -761 389 -749
rect 449 -756 451 -753
rect 459 -756 461 -753
rect 316 -769 318 -765
rect 326 -769 328 -765
rect 387 -774 389 -771
rect 359 -778 361 -775
rect 369 -778 371 -775
rect 415 -776 417 -772
rect 425 -776 427 -772
rect 61 -832 63 -828
rect 71 -832 73 -828
rect 202 -813 204 -809
rect 274 -813 276 -795
rect 284 -813 286 -795
rect 496 -761 498 -758
rect 601 -752 604 -750
rect 644 -752 662 -750
rect 672 -752 675 -750
rect 557 -777 559 -759
rect 567 -777 569 -759
rect 810 -760 812 -757
rect 820 -760 822 -757
rect 860 -758 862 -755
rect 870 -758 872 -755
rect 601 -762 604 -760
rect 644 -762 662 -760
rect 672 -762 675 -760
rect 496 -793 498 -781
rect 161 -825 163 -822
rect 171 -825 173 -822
rect 223 -823 225 -819
rect 233 -823 235 -819
rect 415 -814 417 -796
rect 425 -814 427 -796
rect 449 -814 451 -796
rect 459 -814 461 -796
rect 514 -797 516 -779
rect 524 -797 526 -779
rect 776 -780 778 -776
rect 786 -780 788 -776
rect 599 -787 601 -784
rect 609 -787 611 -784
rect 496 -806 498 -803
rect 557 -801 559 -797
rect 567 -801 569 -797
rect 514 -810 516 -807
rect 524 -810 526 -807
rect 274 -826 276 -823
rect 284 -826 286 -823
rect 127 -836 129 -832
rect 137 -836 139 -832
rect 449 -827 451 -824
rect 459 -827 461 -824
rect 650 -793 652 -789
rect 660 -793 662 -789
rect 681 -799 683 -795
rect 415 -838 417 -834
rect 425 -838 427 -834
rect -144 -855 -142 -843
rect -135 -855 -133 -852
rect 12 -855 14 -852
rect 21 -855 23 -843
rect 599 -845 601 -827
rect 609 -845 611 -827
rect 650 -831 652 -813
rect 660 -831 662 -813
rect 897 -763 899 -759
rect 907 -763 909 -759
rect 987 -763 989 -760
rect 997 -763 999 -760
rect 928 -769 930 -765
rect 776 -818 778 -800
rect 786 -818 788 -800
rect 810 -818 812 -800
rect 820 -818 822 -800
rect 860 -816 862 -798
rect 870 -816 872 -798
rect 897 -801 899 -783
rect 907 -801 909 -783
rect 969 -785 971 -782
rect 928 -801 930 -789
rect 681 -831 683 -819
rect -113 -874 -109 -872
rect -89 -874 -77 -872
rect -67 -874 -63 -872
rect -58 -874 -54 -872
rect -44 -874 -32 -872
rect -12 -874 -8 -872
rect -144 -881 -142 -875
rect -144 -888 -142 -884
rect -135 -888 -133 -875
rect 69 -861 71 -849
rect 78 -861 80 -858
rect 225 -861 227 -858
rect 234 -861 236 -849
rect 12 -888 14 -875
rect 21 -881 23 -875
rect 100 -880 104 -878
rect 124 -880 136 -878
rect 146 -880 150 -878
rect 155 -880 159 -878
rect 169 -880 181 -878
rect 201 -880 205 -878
rect 21 -888 23 -884
rect 69 -887 71 -881
rect 69 -894 71 -890
rect 78 -894 80 -881
rect 357 -863 359 -851
rect 366 -863 368 -860
rect 513 -863 515 -860
rect 522 -863 524 -851
rect 1087 -773 1089 -770
rect 1097 -773 1099 -770
rect 1021 -783 1023 -779
rect 1031 -783 1033 -779
rect 1052 -789 1054 -785
rect 928 -815 930 -811
rect 969 -817 971 -805
rect 897 -825 899 -821
rect 907 -825 909 -821
rect 810 -831 812 -828
rect 820 -831 822 -828
rect 860 -829 862 -826
rect 870 -829 872 -826
rect 987 -821 989 -803
rect 997 -821 999 -803
rect 1021 -821 1023 -803
rect 1031 -821 1033 -803
rect 1052 -821 1054 -809
rect 1115 -795 1117 -792
rect 1146 -795 1148 -791
rect 1156 -795 1158 -791
rect 969 -830 971 -827
rect 987 -834 989 -831
rect 997 -834 999 -831
rect 681 -845 683 -841
rect 776 -842 778 -838
rect 786 -842 788 -838
rect 1087 -831 1089 -813
rect 1097 -831 1099 -813
rect 1115 -827 1117 -815
rect 1052 -835 1054 -831
rect 1146 -833 1148 -815
rect 1156 -833 1158 -815
rect 1115 -840 1117 -837
rect 1021 -845 1023 -841
rect 1031 -845 1033 -841
rect 1087 -844 1089 -841
rect 1097 -844 1099 -841
rect 650 -855 652 -851
rect 660 -855 662 -851
rect 599 -858 601 -855
rect 609 -858 611 -855
rect 225 -894 227 -881
rect 234 -887 236 -881
rect 388 -882 392 -880
rect 412 -882 424 -880
rect 434 -882 438 -880
rect 443 -882 447 -880
rect 457 -882 469 -880
rect 489 -882 493 -880
rect 357 -889 359 -883
rect 234 -894 236 -890
rect -144 -900 -142 -898
rect -144 -904 -143 -900
rect -135 -901 -133 -898
rect 12 -901 14 -898
rect 21 -900 23 -898
rect 22 -904 23 -900
rect 357 -896 359 -892
rect 366 -896 368 -883
rect 718 -867 720 -855
rect 727 -867 729 -864
rect 874 -867 876 -864
rect 883 -867 885 -855
rect 1146 -857 1148 -853
rect 1156 -857 1158 -853
rect 513 -896 515 -883
rect 522 -889 524 -883
rect 749 -886 753 -884
rect 773 -886 785 -884
rect 795 -886 799 -884
rect 804 -886 808 -884
rect 818 -886 830 -884
rect 850 -886 854 -884
rect 522 -896 524 -892
rect 718 -893 720 -887
rect -144 -905 -142 -904
rect 21 -905 23 -904
rect 69 -906 71 -904
rect 69 -910 70 -906
rect 78 -907 80 -904
rect 225 -907 227 -904
rect 234 -906 236 -904
rect 718 -900 720 -896
rect 727 -900 729 -887
rect 1060 -872 1063 -870
rect 1103 -872 1121 -870
rect 1131 -872 1134 -870
rect 950 -877 954 -875
rect 974 -877 992 -875
rect 1012 -877 1016 -875
rect 1060 -882 1063 -880
rect 1103 -882 1121 -880
rect 1131 -882 1134 -880
rect 950 -887 954 -885
rect 974 -887 992 -885
rect 1012 -887 1016 -885
rect 874 -900 876 -887
rect 883 -893 885 -887
rect 883 -900 885 -896
rect 235 -910 236 -906
rect 69 -911 71 -910
rect 234 -911 236 -910
rect 357 -908 359 -906
rect 357 -912 358 -908
rect 366 -909 368 -906
rect 513 -909 515 -906
rect 522 -908 524 -906
rect 523 -912 524 -908
rect 357 -913 359 -912
rect 522 -913 524 -912
rect 718 -912 720 -910
rect 718 -916 719 -912
rect 727 -913 729 -910
rect 874 -913 876 -910
rect 883 -912 885 -910
rect 950 -911 954 -909
rect 974 -911 992 -909
rect 1012 -911 1016 -909
rect 884 -916 885 -912
rect 718 -917 720 -916
rect 883 -917 885 -916
rect 950 -921 954 -919
rect 974 -921 992 -919
rect 1012 -921 1016 -919
<< polycontact >>
rect 228 -706 232 -702
rect 230 -724 234 -720
rect 224 -734 228 -730
rect 312 -738 316 -734
rect 322 -744 326 -740
rect -16 -779 -12 -775
rect -84 -805 -80 -801
rect -74 -799 -70 -795
rect -56 -805 -52 -801
rect -46 -799 -42 -795
rect 8 -805 12 -801
rect 18 -799 22 -795
rect 36 -801 40 -797
rect 57 -801 61 -797
rect 67 -807 71 -803
rect 129 -811 133 -807
rect 139 -805 143 -801
rect 157 -811 161 -807
rect 167 -805 171 -801
rect 204 -798 208 -794
rect 225 -798 229 -794
rect 235 -792 239 -788
rect 355 -764 359 -760
rect 365 -758 369 -754
rect 653 -738 657 -734
rect 383 -760 387 -756
rect 276 -806 280 -802
rect 559 -776 563 -772
rect 651 -756 655 -752
rect 569 -770 573 -766
rect 657 -766 661 -762
rect 498 -792 502 -788
rect 286 -812 290 -808
rect 417 -813 421 -809
rect 427 -807 431 -803
rect 445 -813 449 -809
rect 455 -807 459 -803
rect 516 -790 520 -786
rect 526 -796 530 -792
rect 646 -824 650 -820
rect -142 -848 -138 -844
rect 17 -848 21 -844
rect 595 -844 599 -840
rect 605 -838 609 -834
rect 656 -830 660 -826
rect 893 -794 897 -790
rect 778 -817 782 -813
rect 788 -811 792 -807
rect 806 -817 810 -813
rect 816 -811 820 -807
rect 856 -815 860 -811
rect 866 -809 870 -805
rect 903 -800 907 -796
rect 924 -800 928 -796
rect 677 -830 681 -826
rect -82 -872 -78 -868
rect -43 -872 -39 -868
rect 71 -854 75 -850
rect 230 -854 234 -850
rect -133 -886 -129 -882
rect 8 -886 12 -882
rect 131 -878 135 -874
rect 170 -878 174 -874
rect 359 -856 363 -852
rect 518 -856 522 -852
rect 971 -816 975 -812
rect 989 -814 993 -810
rect 1017 -813 1021 -809
rect 999 -820 1003 -816
rect 1027 -820 1031 -816
rect 1048 -820 1052 -816
rect 1083 -830 1087 -826
rect 1093 -824 1097 -820
rect 1111 -826 1115 -822
rect 1142 -825 1146 -821
rect 1152 -832 1156 -828
rect 80 -892 84 -888
rect 221 -892 225 -888
rect 419 -880 423 -876
rect 458 -880 462 -876
rect -143 -904 -139 -900
rect 18 -904 22 -900
rect 720 -860 724 -856
rect 879 -860 883 -856
rect 368 -894 372 -890
rect 509 -894 513 -890
rect 780 -884 784 -880
rect 819 -884 823 -880
rect 70 -910 74 -906
rect 1116 -870 1120 -866
rect 981 -875 985 -871
rect 987 -885 991 -881
rect 1110 -880 1114 -876
rect 729 -898 733 -894
rect 870 -898 874 -894
rect 231 -910 235 -906
rect 358 -912 362 -908
rect 519 -912 523 -908
rect 981 -909 985 -905
rect 719 -916 723 -912
rect 880 -916 884 -912
rect 987 -919 991 -915
<< metal1 >>
rect 229 -691 269 -688
rect 229 -695 232 -691
rect 227 -698 239 -695
rect 266 -697 269 -691
rect 266 -700 297 -697
rect 310 -700 385 -697
rect 206 -707 217 -704
rect 206 -713 209 -707
rect 229 -713 232 -706
rect 259 -707 286 -704
rect 206 -716 213 -713
rect 206 -731 209 -716
rect 224 -716 241 -713
rect 224 -722 227 -716
rect 223 -725 227 -722
rect -66 -739 -63 -738
rect 209 -735 213 -732
rect -58 -739 38 -738
rect 224 -739 228 -734
rect -66 -741 38 -739
rect -66 -758 -63 -741
rect -57 -748 -54 -741
rect -17 -748 -14 -741
rect 7 -748 10 -741
rect -97 -761 -63 -758
rect 35 -760 38 -741
rect 147 -745 150 -744
rect 231 -741 234 -724
rect 288 -732 291 -709
rect 281 -735 291 -732
rect 155 -745 212 -744
rect 147 -747 212 -745
rect 288 -745 291 -735
rect 294 -734 297 -700
rect 311 -707 314 -700
rect 329 -707 333 -700
rect 354 -707 357 -700
rect 382 -719 385 -700
rect 382 -722 405 -719
rect 321 -728 324 -727
rect 321 -731 333 -728
rect 294 -737 312 -734
rect 330 -740 333 -731
rect 382 -729 385 -722
rect 309 -744 322 -741
rect 330 -743 351 -740
rect 402 -741 405 -722
rect 616 -723 656 -720
rect 500 -732 575 -729
rect 616 -729 619 -723
rect 653 -727 656 -723
rect 588 -732 619 -729
rect 646 -730 658 -727
rect 402 -742 443 -741
rect 330 -745 333 -743
rect -91 -768 -87 -761
rect -72 -768 -69 -761
rect 35 -763 84 -760
rect -8 -775 -5 -768
rect 35 -770 38 -763
rect 56 -770 59 -763
rect 74 -770 78 -763
rect 147 -764 150 -747
rect 156 -754 159 -747
rect 209 -751 212 -747
rect 243 -748 291 -745
rect 243 -751 246 -748
rect 206 -754 246 -751
rect 116 -767 150 -764
rect 206 -767 209 -754
rect 218 -761 222 -754
rect 237 -761 240 -754
rect 288 -755 291 -748
rect 348 -754 351 -743
rect 402 -744 438 -742
rect 348 -757 365 -754
rect 373 -756 376 -747
rect 391 -756 394 -749
rect 435 -747 438 -744
rect 443 -747 472 -746
rect 435 -749 472 -747
rect 373 -759 383 -756
rect 351 -763 355 -760
rect 373 -761 376 -759
rect 391 -759 401 -756
rect 391 -761 394 -759
rect 364 -764 376 -761
rect 364 -765 367 -764
rect 122 -774 126 -767
rect 141 -774 144 -767
rect 311 -770 314 -765
rect 435 -766 438 -749
rect 444 -756 447 -749
rect 500 -761 503 -732
rect 528 -739 531 -732
rect 552 -739 556 -732
rect 571 -739 574 -732
rect 561 -760 564 -759
rect 552 -763 564 -760
rect -23 -778 -16 -775
rect -82 -789 -79 -788
rect -91 -792 -79 -789
rect -91 -801 -88 -792
rect -70 -798 -46 -795
rect -38 -797 -35 -788
rect -38 -800 -32 -797
rect -110 -804 -88 -801
rect -91 -806 -88 -804
rect -80 -805 -56 -802
rect -38 -802 -35 -800
rect -47 -805 -35 -802
rect -23 -802 -20 -778
rect -8 -778 3 -775
rect 302 -773 350 -770
rect 404 -769 438 -766
rect -8 -780 -5 -778
rect -17 -795 -14 -790
rect 0 -795 3 -778
rect 227 -782 230 -781
rect -17 -798 -4 -795
rect 0 -798 18 -795
rect -23 -805 -11 -802
rect -65 -806 -60 -805
rect -47 -806 -44 -805
rect -98 -830 -95 -813
rect -57 -820 -54 -816
rect -38 -819 -35 -816
rect -110 -833 -95 -830
rect -72 -831 -69 -826
rect -66 -823 -38 -820
rect -66 -831 -63 -823
rect -110 -845 -107 -833
rect -72 -834 -63 -831
rect -138 -848 -107 -845
rect -119 -855 -116 -848
rect -128 -858 -79 -855
rect -62 -858 -59 -842
rect -148 -882 -145 -875
rect -82 -868 -79 -858
rect -64 -862 -57 -858
rect -49 -867 -46 -823
rect -14 -826 -11 -805
rect -7 -818 -4 -798
rect 26 -797 29 -788
rect 218 -785 230 -782
rect 44 -797 47 -790
rect 66 -791 69 -790
rect 66 -794 78 -791
rect 26 -800 36 -797
rect 5 -804 8 -801
rect 26 -802 29 -800
rect 44 -800 57 -797
rect 44 -802 47 -800
rect 17 -805 29 -802
rect 17 -806 20 -805
rect 75 -803 78 -794
rect 197 -794 200 -787
rect 218 -794 221 -785
rect 256 -788 259 -782
rect 239 -791 266 -788
rect 131 -795 134 -794
rect 122 -798 134 -795
rect 55 -807 67 -804
rect 75 -806 84 -803
rect 75 -808 78 -806
rect 7 -820 10 -816
rect 26 -820 29 -816
rect 35 -819 38 -812
rect -3 -823 34 -820
rect 81 -824 84 -806
rect -14 -829 1 -826
rect -2 -835 1 -829
rect 81 -827 97 -824
rect 56 -832 59 -828
rect 108 -830 111 -800
rect 122 -807 125 -798
rect 143 -804 167 -801
rect 175 -803 178 -794
rect 194 -797 200 -794
rect 197 -799 200 -797
rect 208 -797 221 -794
rect 218 -799 221 -797
rect 229 -798 248 -795
rect 175 -806 187 -803
rect 263 -804 266 -791
rect 269 -804 272 -795
rect 119 -810 125 -807
rect 122 -812 125 -810
rect 133 -811 157 -808
rect 175 -808 178 -806
rect 166 -811 178 -808
rect 184 -809 187 -806
rect 263 -807 272 -804
rect 280 -805 293 -802
rect 148 -812 153 -811
rect 166 -812 169 -811
rect 2 -839 42 -836
rect 91 -833 111 -830
rect 60 -836 81 -833
rect 91 -841 94 -833
rect 115 -836 118 -819
rect 156 -826 159 -822
rect 175 -824 178 -822
rect 206 -823 209 -809
rect 269 -809 272 -807
rect 269 -812 281 -809
rect 290 -811 298 -808
rect 278 -813 281 -812
rect 175 -826 205 -824
rect 147 -827 205 -826
rect 103 -839 118 -836
rect 141 -837 144 -832
rect 147 -829 178 -827
rect 237 -824 240 -819
rect 210 -827 246 -824
rect 269 -827 272 -823
rect 288 -827 291 -823
rect 302 -827 305 -773
rect 347 -779 350 -773
rect 354 -779 357 -775
rect 373 -779 376 -775
rect 382 -779 385 -771
rect 347 -782 385 -779
rect 410 -776 414 -769
rect 429 -776 432 -769
rect 552 -772 555 -763
rect 588 -766 591 -732
rect 573 -769 591 -766
rect 599 -739 626 -736
rect 594 -764 597 -741
rect 653 -745 656 -738
rect 668 -739 679 -736
rect 676 -745 679 -739
rect 644 -748 661 -745
rect 658 -754 661 -748
rect 672 -748 679 -745
rect 594 -767 604 -764
rect 534 -775 555 -772
rect 147 -837 150 -829
rect -16 -847 -15 -842
rect -10 -845 -9 -842
rect -10 -847 17 -845
rect -16 -848 17 -847
rect -16 -849 -9 -848
rect -5 -855 -2 -848
rect 103 -851 106 -839
rect 141 -840 150 -837
rect 75 -854 106 -851
rect -67 -870 -54 -867
rect -47 -871 -46 -867
rect -42 -858 7 -855
rect -42 -868 -39 -858
rect 94 -861 97 -854
rect 85 -864 134 -861
rect 151 -864 154 -848
rect -140 -876 -137 -873
rect -89 -879 -77 -876
rect -44 -879 -32 -876
rect 16 -876 19 -873
rect -157 -884 -145 -882
rect -152 -885 -145 -884
rect -148 -888 -145 -885
rect -140 -888 -137 -881
rect -129 -886 -123 -883
rect -82 -887 -79 -879
rect -112 -890 -79 -887
rect -42 -887 -39 -879
rect 2 -886 8 -883
rect -42 -890 -9 -887
rect 16 -888 19 -881
rect -112 -893 -109 -890
rect -125 -895 -109 -893
rect -128 -896 -109 -895
rect -12 -893 -9 -890
rect 24 -882 27 -875
rect 24 -884 36 -882
rect 24 -885 31 -884
rect 24 -888 27 -885
rect 65 -888 68 -881
rect 131 -874 134 -864
rect 149 -868 156 -864
rect 164 -873 167 -829
rect 242 -830 305 -827
rect 382 -824 385 -782
rect 491 -788 494 -781
rect 509 -788 512 -779
rect 534 -786 537 -775
rect 552 -777 555 -775
rect 563 -776 577 -773
rect 594 -777 597 -767
rect 651 -773 654 -756
rect 658 -757 662 -754
rect 676 -763 679 -748
rect 796 -751 799 -750
rect 842 -750 889 -748
rect 804 -751 889 -750
rect 796 -753 845 -751
rect 657 -769 661 -766
rect 672 -767 676 -764
rect 594 -780 642 -777
rect 796 -770 799 -753
rect 805 -760 808 -753
rect 855 -758 858 -751
rect 886 -753 889 -751
rect 886 -756 1014 -753
rect 892 -763 895 -756
rect 910 -763 914 -756
rect 760 -773 799 -770
rect 923 -769 926 -756
rect 482 -791 494 -788
rect 419 -797 422 -796
rect 410 -800 422 -797
rect 396 -832 399 -802
rect 410 -807 413 -800
rect 431 -806 455 -803
rect 463 -805 466 -796
rect 482 -799 485 -791
rect 491 -793 494 -791
rect 502 -791 512 -788
rect 520 -789 537 -786
rect 594 -787 597 -780
rect 639 -783 642 -780
rect 760 -783 763 -773
rect 639 -786 763 -783
rect 771 -780 775 -773
rect 790 -780 793 -773
rect 973 -775 976 -756
rect 1001 -763 1004 -756
rect 962 -778 976 -775
rect 1011 -773 1014 -756
rect 1047 -766 1113 -763
rect 1047 -773 1050 -766
rect 1011 -776 1050 -773
rect 902 -784 905 -783
rect 509 -793 512 -791
rect 509 -796 521 -793
rect 530 -795 534 -792
rect 518 -797 521 -796
rect 645 -793 648 -786
rect 663 -793 667 -786
rect 571 -802 574 -797
rect 676 -799 679 -786
rect 902 -787 914 -784
rect 973 -785 976 -778
rect 891 -794 893 -790
rect 409 -812 413 -807
rect 463 -808 475 -805
rect 410 -814 413 -812
rect 421 -813 445 -810
rect 463 -810 466 -808
rect 454 -813 466 -810
rect 472 -810 475 -808
rect 436 -814 441 -813
rect 454 -814 457 -813
rect 500 -811 503 -803
rect 509 -811 512 -807
rect 528 -811 531 -807
rect 535 -805 583 -802
rect 911 -796 914 -787
rect 1016 -783 1019 -776
rect 1034 -783 1038 -776
rect 1047 -789 1050 -776
rect 1082 -773 1085 -766
rect 1110 -785 1113 -766
rect 1110 -788 1169 -785
rect 932 -796 935 -789
rect 1110 -795 1113 -788
rect 1141 -795 1144 -788
rect 1159 -795 1163 -788
rect 780 -801 783 -800
rect 535 -811 538 -805
rect 500 -814 538 -811
rect 379 -835 399 -832
rect 211 -841 214 -839
rect 379 -843 382 -835
rect 403 -838 406 -821
rect 444 -828 447 -824
rect 463 -826 466 -824
rect 463 -828 464 -826
rect 391 -841 406 -838
rect 429 -839 432 -834
rect 435 -831 464 -828
rect 435 -839 438 -831
rect 197 -853 198 -848
rect 203 -851 204 -848
rect 203 -853 230 -851
rect 197 -854 230 -853
rect 197 -855 204 -854
rect 208 -861 211 -854
rect 391 -853 394 -841
rect 429 -842 438 -839
rect 363 -856 394 -853
rect 146 -876 159 -873
rect 166 -877 167 -873
rect 171 -864 220 -861
rect 171 -874 174 -864
rect 382 -863 385 -856
rect 373 -866 422 -863
rect 439 -866 442 -850
rect 73 -882 76 -879
rect 124 -885 136 -882
rect 169 -885 181 -882
rect 229 -882 232 -879
rect 56 -890 68 -888
rect -12 -895 4 -893
rect -12 -896 7 -895
rect -128 -898 -122 -896
rect -125 -901 -122 -898
rect -139 -904 -122 -901
rect 1 -898 7 -896
rect 61 -891 68 -890
rect 65 -894 68 -891
rect 73 -894 76 -887
rect 84 -892 90 -889
rect 131 -893 134 -885
rect 101 -896 134 -893
rect 171 -893 174 -885
rect 215 -892 221 -889
rect 171 -896 204 -893
rect 229 -894 232 -887
rect 1 -901 4 -898
rect 101 -899 104 -896
rect 1 -904 18 -901
rect 88 -901 104 -899
rect 85 -902 104 -901
rect 201 -899 204 -896
rect 237 -888 240 -881
rect 237 -890 249 -888
rect 353 -890 356 -883
rect 419 -876 422 -866
rect 437 -870 444 -866
rect 452 -875 455 -831
rect 485 -855 486 -850
rect 491 -853 492 -850
rect 491 -855 518 -853
rect 485 -856 518 -855
rect 485 -857 492 -856
rect 496 -863 499 -856
rect 580 -859 583 -805
rect 771 -804 783 -801
rect 655 -814 658 -813
rect 655 -817 667 -814
rect 619 -823 646 -820
rect 592 -837 605 -834
rect 613 -836 616 -827
rect 619 -836 622 -823
rect 664 -826 667 -817
rect 685 -826 688 -819
rect 643 -830 656 -827
rect 664 -829 677 -826
rect 664 -831 667 -829
rect 685 -829 691 -826
rect 685 -831 688 -829
rect 757 -836 760 -806
rect 771 -811 774 -804
rect 792 -810 816 -807
rect 824 -809 827 -800
rect 835 -808 866 -805
rect 835 -809 838 -808
rect 874 -807 877 -798
rect 886 -800 903 -797
rect 911 -799 924 -796
rect 886 -807 889 -800
rect 911 -801 914 -799
rect 932 -799 944 -796
rect 932 -801 935 -799
rect 770 -816 774 -811
rect 824 -812 838 -809
rect 874 -810 889 -807
rect 771 -818 774 -816
rect 782 -817 806 -814
rect 824 -814 827 -812
rect 815 -817 827 -814
rect 797 -818 802 -817
rect 815 -818 818 -817
rect 831 -819 834 -812
rect 852 -814 856 -811
rect 874 -812 877 -810
rect 865 -815 877 -812
rect 941 -810 944 -799
rect 865 -816 868 -815
rect 613 -839 622 -836
rect 587 -843 595 -840
rect 613 -841 616 -839
rect 604 -844 616 -841
rect 740 -839 760 -836
rect 604 -845 607 -844
rect 594 -859 597 -855
rect 613 -859 616 -855
rect 645 -856 648 -851
rect 676 -855 679 -841
rect 740 -847 743 -839
rect 764 -842 767 -825
rect 805 -832 808 -828
rect 824 -830 827 -828
rect 892 -826 895 -821
rect 923 -826 926 -811
rect 964 -812 967 -805
rect 982 -812 985 -803
rect 1026 -804 1029 -803
rect 1026 -807 1038 -804
rect 957 -815 967 -812
rect 964 -817 967 -815
rect 975 -815 985 -812
rect 993 -813 1017 -810
rect 982 -817 985 -815
rect 1035 -816 1038 -807
rect 1056 -816 1059 -809
rect 982 -820 994 -817
rect 1003 -819 1027 -816
rect 1035 -819 1048 -816
rect 991 -821 994 -820
rect 1035 -821 1038 -819
rect 1056 -821 1063 -816
rect 855 -830 858 -826
rect 874 -830 877 -826
rect 886 -829 926 -826
rect 1059 -825 1063 -821
rect 1080 -823 1093 -820
rect 1101 -822 1104 -813
rect 1119 -822 1122 -815
rect 1151 -816 1154 -815
rect 1151 -819 1163 -816
rect 886 -830 889 -829
rect 824 -832 889 -830
rect 796 -833 889 -832
rect 752 -845 767 -842
rect 790 -843 793 -838
rect 796 -835 827 -833
rect 923 -835 926 -829
rect 973 -835 976 -827
rect 982 -835 985 -831
rect 1001 -835 1004 -831
rect 796 -843 799 -835
rect 639 -859 675 -856
rect 580 -862 643 -859
rect 752 -857 755 -845
rect 790 -846 799 -843
rect 724 -860 755 -857
rect 434 -878 447 -875
rect 454 -879 455 -875
rect 459 -866 508 -863
rect 459 -876 462 -866
rect 743 -867 746 -860
rect 734 -870 783 -867
rect 800 -870 803 -854
rect 361 -884 364 -881
rect 412 -887 424 -884
rect 457 -887 469 -884
rect 517 -884 520 -881
rect 237 -891 244 -890
rect 237 -894 240 -891
rect 344 -892 356 -890
rect 349 -893 356 -892
rect 353 -896 356 -893
rect 201 -901 217 -899
rect 361 -896 364 -889
rect 372 -894 378 -891
rect 419 -895 422 -887
rect 389 -898 422 -895
rect 459 -895 462 -887
rect 503 -894 509 -891
rect 459 -898 492 -895
rect 517 -896 520 -889
rect 201 -902 220 -901
rect 85 -904 91 -902
rect 88 -907 91 -904
rect 74 -910 91 -907
rect 214 -904 220 -902
rect 389 -901 392 -898
rect 214 -907 217 -904
rect 376 -903 392 -901
rect 373 -904 392 -903
rect 489 -901 492 -898
rect 525 -890 528 -883
rect 525 -892 537 -890
rect 525 -893 532 -892
rect 525 -896 528 -893
rect 714 -894 717 -887
rect 780 -880 783 -870
rect 798 -874 805 -870
rect 813 -879 816 -835
rect 923 -838 1012 -835
rect 860 -848 863 -844
rect 1009 -846 1012 -838
rect 1016 -846 1019 -841
rect 1047 -845 1050 -831
rect 1060 -834 1063 -825
rect 1101 -825 1111 -822
rect 1075 -828 1083 -827
rect 1080 -830 1083 -828
rect 1101 -827 1104 -825
rect 1119 -825 1142 -822
rect 1119 -827 1122 -825
rect 1092 -830 1104 -827
rect 1092 -831 1095 -830
rect 1160 -828 1163 -819
rect 1061 -839 1063 -834
rect 1141 -832 1152 -829
rect 1160 -831 1173 -828
rect 1160 -833 1163 -831
rect 1082 -845 1085 -841
rect 1101 -845 1104 -841
rect 1110 -845 1113 -837
rect 1047 -846 1138 -845
rect 1009 -848 1138 -846
rect 1009 -849 1050 -848
rect 846 -859 847 -854
rect 852 -857 853 -854
rect 852 -859 879 -857
rect 846 -860 879 -859
rect 846 -861 853 -860
rect 857 -867 860 -860
rect 795 -882 808 -879
rect 815 -883 816 -879
rect 820 -870 869 -867
rect 820 -880 823 -870
rect 944 -870 947 -864
rect 944 -873 954 -870
rect 722 -888 725 -885
rect 773 -891 785 -888
rect 818 -891 830 -888
rect 878 -888 881 -885
rect 705 -896 717 -894
rect 710 -897 717 -896
rect 714 -900 717 -897
rect 489 -903 505 -901
rect 489 -904 508 -903
rect 373 -906 379 -904
rect 214 -910 231 -907
rect 376 -909 379 -906
rect 362 -912 379 -909
rect 502 -906 508 -904
rect 722 -900 725 -893
rect 733 -898 739 -895
rect 780 -899 783 -891
rect 750 -902 783 -899
rect 820 -899 823 -891
rect 864 -898 870 -895
rect 820 -902 853 -899
rect 878 -900 881 -893
rect 750 -905 753 -902
rect 502 -909 505 -906
rect 502 -912 519 -909
rect 737 -907 753 -905
rect 734 -908 753 -907
rect 850 -905 853 -902
rect 886 -894 889 -887
rect 944 -888 947 -873
rect 981 -871 984 -862
rect 988 -864 991 -856
rect 988 -869 989 -864
rect 974 -883 978 -880
rect 988 -881 991 -869
rect 1017 -870 1020 -849
rect 1012 -873 1020 -870
rect 944 -892 954 -888
rect 975 -889 978 -883
rect 975 -892 992 -889
rect 886 -896 898 -894
rect 886 -897 893 -896
rect 886 -900 889 -897
rect 944 -904 947 -892
rect 850 -907 866 -905
rect 850 -908 869 -907
rect 734 -910 740 -908
rect 737 -913 740 -910
rect 723 -916 740 -913
rect 863 -910 869 -908
rect 944 -907 954 -904
rect 863 -913 866 -910
rect 863 -916 880 -913
rect 944 -922 947 -907
rect 981 -905 985 -903
rect 974 -917 978 -914
rect 988 -915 991 -892
rect 1017 -904 1020 -873
rect 1053 -865 1056 -863
rect 1053 -868 1063 -865
rect 1053 -893 1056 -868
rect 1110 -876 1113 -851
rect 1135 -858 1138 -848
rect 1170 -851 1173 -831
rect 1141 -858 1144 -853
rect 1135 -861 1166 -858
rect 1116 -866 1119 -861
rect 1135 -865 1138 -861
rect 1131 -868 1138 -865
rect 1117 -878 1121 -875
rect 1117 -884 1120 -878
rect 1103 -887 1120 -884
rect 1135 -884 1138 -868
rect 1131 -887 1138 -884
rect 1112 -898 1115 -887
rect 1046 -901 1115 -898
rect 1012 -907 1020 -904
rect 944 -926 954 -922
rect 975 -923 978 -917
rect 975 -926 992 -923
rect 944 -932 947 -926
rect 987 -932 990 -926
rect 1017 -929 1020 -907
<< m2contact >>
rect 305 -700 310 -695
rect 286 -709 291 -704
rect 222 -744 227 -739
rect 231 -746 236 -741
rect 575 -732 580 -727
rect -106 -794 -100 -789
rect -115 -805 -110 -800
rect -65 -795 -60 -790
rect -32 -801 -27 -796
rect -99 -813 -94 -808
rect -65 -811 -60 -806
rect -123 -840 -118 -835
rect -69 -863 -64 -858
rect -57 -863 -52 -858
rect -38 -824 -33 -819
rect 0 -806 5 -801
rect 108 -800 113 -795
rect 50 -809 55 -804
rect -8 -823 -3 -818
rect 34 -824 39 -819
rect 97 -827 102 -822
rect 114 -810 119 -805
rect 148 -801 153 -796
rect 189 -799 194 -794
rect 293 -805 298 -800
rect 114 -819 119 -814
rect 148 -817 153 -812
rect 184 -814 189 -809
rect -3 -840 2 -835
rect 55 -837 60 -832
rect 294 -816 299 -811
rect 594 -741 599 -736
rect 90 -846 95 -841
rect -141 -881 -136 -876
rect 15 -881 20 -876
rect 144 -869 149 -864
rect 156 -869 161 -864
rect 577 -777 582 -772
rect 649 -778 654 -773
rect 396 -802 401 -797
rect 382 -829 387 -824
rect 436 -803 441 -798
rect 886 -794 891 -789
rect 403 -812 409 -807
rect 402 -821 407 -816
rect 436 -819 441 -814
rect 472 -815 477 -810
rect 210 -846 215 -841
rect 464 -831 469 -826
rect 378 -848 383 -843
rect 72 -887 77 -882
rect 228 -887 233 -882
rect 432 -871 437 -866
rect 444 -871 449 -866
rect 498 -848 503 -843
rect 757 -806 762 -801
rect 587 -837 592 -832
rect 691 -831 696 -826
rect 797 -807 802 -802
rect 765 -816 770 -811
rect 763 -825 768 -820
rect 797 -823 802 -818
rect 847 -816 852 -811
rect 830 -824 835 -819
rect 586 -848 591 -843
rect 1075 -824 1080 -819
rect 739 -852 744 -847
rect 360 -889 365 -884
rect 516 -889 521 -884
rect 793 -875 798 -870
rect 805 -875 810 -870
rect 1075 -833 1080 -828
rect 1056 -839 1061 -834
rect 1136 -833 1141 -828
rect 859 -853 864 -848
rect 943 -864 948 -859
rect 721 -893 726 -888
rect 877 -893 882 -888
rect 989 -869 994 -864
rect 1105 -856 1110 -851
rect 980 -903 985 -898
rect 1116 -861 1121 -856
rect 1170 -856 1175 -851
rect 1041 -901 1046 -896
<< pdm12contact >>
rect -109 -871 -104 -866
rect -17 -871 -12 -866
rect 104 -877 109 -872
rect 196 -877 201 -872
rect 392 -879 397 -874
rect 484 -879 489 -874
rect 753 -883 758 -878
rect 845 -883 850 -878
<< metal2 >>
rect 288 -699 305 -696
rect 288 -704 291 -699
rect 140 -735 163 -732
rect 140 -756 143 -735
rect 160 -741 163 -735
rect 580 -731 597 -728
rect 594 -736 597 -731
rect 160 -744 222 -741
rect 236 -745 298 -742
rect 51 -759 143 -756
rect 51 -781 54 -759
rect 190 -760 249 -757
rect -114 -784 54 -781
rect -114 -800 -111 -784
rect -100 -793 -65 -790
rect -106 -825 -103 -794
rect -31 -802 -27 -801
rect -31 -805 0 -802
rect -94 -811 -65 -808
rect 51 -804 54 -784
rect 100 -806 103 -773
rect 190 -794 193 -760
rect 113 -799 148 -796
rect 295 -800 298 -745
rect 578 -772 581 -762
rect 587 -777 649 -774
rect 577 -783 580 -777
rect 258 -804 293 -801
rect 100 -809 114 -806
rect -33 -823 -8 -820
rect 119 -817 148 -814
rect 258 -810 261 -804
rect 388 -786 580 -783
rect 298 -804 343 -801
rect 189 -813 261 -810
rect 299 -815 317 -811
rect 39 -823 55 -820
rect -114 -828 -103 -825
rect -114 -836 -111 -828
rect -118 -839 -111 -836
rect -161 -877 -158 -849
rect -161 -880 -141 -877
rect -122 -882 -119 -840
rect 52 -836 55 -823
rect 102 -826 120 -823
rect -108 -854 -73 -851
rect -108 -866 -105 -854
rect -76 -859 -73 -854
rect -48 -854 -13 -851
rect -76 -862 -69 -859
rect -48 -859 -45 -854
rect -52 -862 -45 -859
rect -16 -866 -13 -854
rect -2 -882 1 -840
rect 117 -834 120 -826
rect 117 -837 214 -834
rect 211 -841 214 -837
rect 340 -835 343 -804
rect 388 -808 391 -786
rect 401 -801 436 -798
rect 388 -811 403 -808
rect 407 -819 436 -816
rect 473 -818 577 -815
rect 387 -829 464 -826
rect 574 -834 577 -818
rect 587 -832 590 -777
rect 650 -781 841 -778
rect 636 -792 695 -789
rect 692 -826 695 -792
rect 762 -805 797 -802
rect 750 -815 765 -812
rect 750 -832 753 -815
rect 838 -812 841 -781
rect 887 -789 890 -741
rect 838 -815 847 -812
rect 1068 -818 1071 -793
rect 768 -823 797 -820
rect 1068 -819 1078 -818
rect 1068 -821 1075 -819
rect 831 -825 835 -824
rect 831 -828 1068 -825
rect 1065 -829 1068 -828
rect 1065 -832 1075 -829
rect 340 -838 564 -835
rect 574 -837 587 -834
rect 750 -835 920 -832
rect 1132 -832 1136 -829
rect 20 -880 43 -877
rect 40 -906 43 -880
rect 52 -883 55 -855
rect 52 -886 72 -883
rect 91 -888 94 -846
rect 215 -845 282 -842
rect 105 -860 140 -857
rect 105 -872 108 -860
rect 137 -865 140 -860
rect 165 -860 200 -857
rect 137 -868 144 -865
rect 165 -865 168 -860
rect 161 -868 168 -865
rect 197 -872 200 -860
rect 211 -888 214 -846
rect 233 -886 256 -883
rect 253 -912 256 -886
rect 340 -885 343 -857
rect 340 -888 360 -885
rect 379 -890 382 -848
rect 561 -844 564 -838
rect 561 -847 586 -844
rect 393 -862 428 -859
rect 393 -874 396 -862
rect 425 -867 428 -862
rect 453 -862 488 -859
rect 425 -870 432 -867
rect 453 -867 456 -862
rect 449 -870 456 -867
rect 485 -874 488 -862
rect 499 -890 502 -848
rect 521 -888 544 -885
rect 541 -914 544 -888
rect 701 -889 704 -861
rect 701 -892 721 -889
rect 740 -894 743 -852
rect 917 -850 920 -835
rect 917 -853 927 -850
rect 754 -866 789 -863
rect 754 -878 757 -866
rect 786 -871 789 -866
rect 814 -866 849 -863
rect 786 -874 793 -871
rect 814 -871 817 -866
rect 810 -874 817 -871
rect 846 -878 849 -866
rect 860 -894 863 -853
rect 1057 -850 1060 -839
rect 1057 -851 1110 -850
rect 1057 -853 1105 -851
rect 1116 -855 1170 -852
rect 1116 -856 1121 -855
rect 948 -863 952 -860
rect 1040 -862 1051 -859
rect 994 -869 1030 -866
rect 1027 -884 1030 -869
rect 882 -892 905 -889
rect 902 -918 905 -892
rect 981 -898 1041 -897
rect 985 -900 1041 -898
<< m3contact >>
rect 99 -773 104 -768
rect -31 -810 -26 -805
rect 249 -761 254 -756
rect 317 -816 322 -811
rect -162 -849 -157 -844
rect 631 -793 636 -788
rect 51 -855 56 -850
rect 282 -846 287 -841
rect 339 -857 344 -852
rect 700 -861 705 -856
rect 927 -854 932 -849
<< m123contact >>
rect -63 -739 -58 -734
rect 150 -745 155 -740
rect 204 -736 209 -731
rect 304 -745 309 -740
rect 255 -782 260 -777
rect 248 -799 253 -794
rect 438 -747 443 -742
rect 799 -751 804 -746
rect 346 -765 351 -760
rect 676 -768 681 -763
rect -63 -842 -58 -837
rect -15 -847 -10 -842
rect 205 -828 210 -823
rect 534 -797 539 -792
rect 481 -804 486 -799
rect 658 -774 663 -769
rect 638 -831 643 -826
rect 957 -778 962 -773
rect 940 -815 945 -810
rect -157 -889 -152 -884
rect -123 -887 -118 -882
rect -3 -887 2 -882
rect 31 -889 36 -884
rect 150 -848 155 -843
rect 198 -853 203 -848
rect 56 -895 61 -890
rect 90 -893 95 -888
rect 210 -893 215 -888
rect 244 -895 249 -890
rect 438 -850 443 -845
rect 859 -844 864 -839
rect 486 -855 491 -850
rect 675 -860 680 -855
rect 344 -897 349 -892
rect 378 -895 383 -890
rect 498 -895 503 -890
rect 532 -897 537 -892
rect 799 -854 804 -849
rect 847 -859 852 -854
rect 980 -862 985 -857
rect 1051 -863 1056 -858
rect 705 -901 710 -896
rect 739 -899 744 -894
rect 859 -899 864 -894
rect 893 -901 898 -896
<< metal3 >>
rect 195 -727 304 -724
rect 135 -731 168 -728
rect -62 -837 -59 -739
rect 135 -751 138 -731
rect 165 -736 168 -731
rect 195 -736 198 -727
rect 165 -739 198 -736
rect 100 -754 138 -751
rect 100 -767 103 -754
rect 98 -768 105 -767
rect 98 -773 99 -768
rect 104 -773 105 -768
rect 98 -774 105 -773
rect -32 -805 -25 -804
rect -32 -810 -31 -805
rect -26 -810 -25 -805
rect -32 -811 -25 -810
rect -31 -827 -27 -811
rect 93 -827 97 -793
rect -31 -831 97 -827
rect -163 -844 -156 -843
rect -163 -849 -162 -844
rect -157 -846 -156 -844
rect -16 -846 -15 -842
rect -157 -847 -15 -846
rect -10 -847 -9 -842
rect 151 -843 154 -745
rect 205 -823 208 -736
rect 301 -744 304 -727
rect 428 -737 451 -734
rect 305 -749 308 -745
rect 428 -749 431 -737
rect 448 -741 451 -737
rect 448 -744 649 -741
rect 305 -752 431 -749
rect 248 -756 255 -755
rect 248 -761 249 -756
rect 254 -757 255 -756
rect 254 -760 347 -757
rect 254 -761 255 -760
rect 248 -762 255 -761
rect 344 -763 346 -760
rect 255 -777 260 -774
rect -157 -849 -9 -847
rect -163 -850 -156 -849
rect 50 -850 57 -849
rect 50 -855 51 -850
rect 56 -852 57 -850
rect 197 -852 198 -848
rect 56 -853 198 -852
rect 203 -853 204 -848
rect 56 -855 204 -853
rect 50 -856 57 -855
rect 249 -869 252 -799
rect 317 -810 321 -793
rect 316 -811 323 -810
rect 316 -816 317 -811
rect 322 -816 323 -811
rect 316 -817 323 -816
rect 281 -841 288 -840
rect 281 -846 282 -841
rect 287 -844 355 -841
rect 287 -846 288 -844
rect 439 -845 442 -747
rect 646 -769 649 -744
rect 646 -772 658 -769
rect 630 -788 637 -787
rect 630 -789 631 -788
rect 538 -792 631 -789
rect 539 -795 541 -792
rect 630 -793 631 -792
rect 636 -793 637 -788
rect 630 -794 637 -793
rect 482 -822 485 -804
rect 482 -825 498 -822
rect 628 -830 638 -827
rect 281 -847 288 -846
rect 338 -852 345 -851
rect 338 -857 339 -852
rect 344 -854 345 -852
rect 485 -854 486 -850
rect 344 -855 486 -854
rect 491 -855 492 -850
rect 628 -851 631 -830
rect 567 -854 631 -851
rect 677 -855 680 -768
rect 800 -849 803 -751
rect 941 -838 944 -815
rect 958 -831 961 -778
rect 958 -834 972 -831
rect 840 -844 859 -841
rect 941 -841 963 -838
rect 926 -849 933 -848
rect 926 -854 927 -849
rect 932 -852 940 -849
rect 932 -854 933 -852
rect 344 -857 492 -855
rect 338 -858 345 -857
rect 699 -856 706 -855
rect 699 -861 700 -856
rect 705 -858 706 -856
rect 846 -858 847 -854
rect 705 -859 847 -858
rect 852 -859 853 -854
rect 926 -855 933 -854
rect 960 -853 963 -841
rect 969 -840 972 -834
rect 969 -843 1008 -840
rect 1005 -851 1008 -843
rect 960 -856 984 -853
rect 1005 -854 1055 -851
rect 705 -861 853 -859
rect 980 -857 984 -856
rect 699 -862 706 -861
rect 1052 -858 1055 -854
rect 114 -872 252 -869
rect -155 -884 -123 -883
rect -152 -886 -123 -884
rect 2 -884 34 -883
rect 2 -886 31 -884
rect 32 -902 35 -889
rect 58 -890 90 -889
rect 61 -892 90 -890
rect 114 -902 117 -872
rect 215 -890 247 -889
rect 215 -892 244 -890
rect 346 -892 378 -891
rect 349 -894 378 -892
rect 503 -892 535 -891
rect 503 -894 532 -892
rect 707 -896 739 -895
rect 710 -898 739 -896
rect 864 -896 896 -895
rect 864 -898 893 -896
rect 32 -905 117 -902
<< m234contact >>
rect 38 -841 43 -836
rect 886 -741 891 -736
rect 577 -762 582 -757
rect 1067 -793 1072 -788
rect 1127 -833 1132 -828
rect 952 -865 957 -860
rect 1035 -864 1040 -859
rect 1026 -889 1031 -884
<< m4contact >>
rect 93 -793 98 -788
rect 255 -774 260 -769
rect 317 -793 322 -788
rect 355 -844 360 -839
rect 498 -825 503 -820
rect 562 -855 567 -850
rect 835 -845 840 -840
rect 940 -852 945 -847
<< metal4 >>
rect 256 -713 411 -710
rect 256 -769 259 -713
rect 408 -720 411 -713
rect 606 -713 673 -710
rect 606 -720 609 -713
rect 408 -723 609 -720
rect 670 -725 673 -713
rect 670 -728 689 -725
rect 686 -754 689 -728
rect 785 -740 886 -737
rect 785 -754 788 -740
rect 686 -757 788 -754
rect 947 -753 1071 -750
rect 582 -761 632 -758
rect 98 -793 317 -789
rect 629 -805 632 -761
rect 947 -805 950 -753
rect 1068 -788 1071 -753
rect 629 -808 950 -805
rect 503 -824 737 -821
rect 39 -909 42 -841
rect 360 -843 555 -840
rect 552 -852 555 -843
rect 734 -842 737 -824
rect 734 -845 835 -842
rect 552 -855 562 -852
rect 1128 -848 1131 -833
rect 945 -851 1131 -848
rect 957 -863 1035 -860
rect 630 -871 916 -868
rect 630 -893 633 -871
rect 138 -896 633 -893
rect 138 -898 141 -896
rect 110 -901 141 -898
rect 110 -909 113 -901
rect 39 -912 113 -909
rect 913 -913 916 -871
rect 1027 -913 1030 -889
rect 913 -916 1030 -913
<< labels >>
rlabel metal1 -61 -860 -61 -860 3 vdd
rlabel metal1 -61 -868 -61 -868 3 gnd
rlabel metal1 -75 -760 -75 -760 5 vdd
rlabel metal1 -46 -821 -46 -821 1 gnd
rlabel metal1 -56 -740 -56 -739 5 vdd
rlabel metal1 78 -806 84 -803 7 c1
rlabel metal1 71 -835 71 -835 1 gnd
rlabel metal1 62 -762 62 -762 5 vdd
rlabel m2contact 1 -803 5 -802 1 p0_inv
rlabel metal1 45 -799 47 -796 1 temp100
rlabel metal1 8 -740 8 -739 5 vdd
rlabel metal1 18 -821 18 -821 1 gnd
rlabel metal1 -7 -777 -5 -774 1 c0_inv
rlabel metal1 -22 -778 -20 -776 3 c0
rlabel metal1 -16 -797 -16 -797 1 gnd
rlabel metal1 -17 -739 -17 -739 5 vdd
rlabel m2contact -1 -838 0 -838 1 c0
rlabel metal2 41 -906 42 -904 1 s0
rlabel metal2 -160 -879 -156 -877 3 mid_s0
rlabel metal1 -68 -798 -57 -795 1 a0
rlabel metal1 -68 -805 -57 -802 1 b0
rlabel metal1 -97 -804 -91 -801 1 g0_inv
rlabel metal1 -35 -800 -30 -797 1 p0_inv
rlabel m2contact 51 -807 55 -805 1 g0_inv
rlabel metal1 152 -866 152 -866 3 vdd
rlabel metal1 152 -874 152 -874 3 gnd
rlabel metal1 138 -766 138 -766 5 vdd
rlabel metal1 167 -827 167 -827 1 gnd
rlabel metal1 157 -746 157 -745 5 vdd
rlabel metal2 53 -884 53 -884 1 mid_s1
rlabel metal2 254 -912 255 -910 8 s1
rlabel metal1 116 -810 122 -807 1 g1_inv
rlabel metal1 178 -806 183 -803 1 p1_inv
rlabel metal1 145 -804 156 -801 1 a1
rlabel metal1 145 -811 156 -808 1 b1
rlabel metal1 212 -842 214 -839 1 c1
rlabel metal1 290 -747 290 -746 5 vdd
rlabel metal1 280 -828 280 -828 1 gnd
rlabel metal1 291 -805 295 -803 7 p1_inv
rlabel metal1 292 -811 297 -809 7 p0_inv
rlabel metal1 264 -807 268 -805 3 temp101
rlabel metal1 234 -753 234 -753 5 vdd
rlabel metal1 225 -826 225 -826 1 gnd
rlabel metal1 241 -797 245 -796 1 c0
rlabel metal1 197 -796 199 -794 1 temp102
rlabel metal1 208 -724 208 -724 3 gnd
rlabel metal1 289 -734 290 -734 7 vdd
rlabel space 225 -740 228 -737 1 g0_inv
rlabel metal1 230 -698 233 -695 1 temp103
rlabel metal1 317 -699 317 -699 5 vdd
rlabel metal1 326 -772 326 -772 1 gnd
rlabel metal1 333 -743 339 -740 7 temp104
rlabel metal1 355 -699 355 -698 5 vdd
rlabel metal1 365 -780 365 -780 1 gnd
rlabel metal1 392 -758 394 -756 1 c2
rlabel m123contact 305 -743 305 -743 1 g1_inv
rlabel metal1 440 -868 440 -868 3 vdd
rlabel metal1 440 -876 440 -876 3 gnd
rlabel metal1 426 -768 426 -768 5 vdd
rlabel metal1 455 -829 455 -829 1 gnd
rlabel metal1 445 -748 445 -747 5 vdd
rlabel metal2 342 -887 343 -885 1 mid_s2
rlabel metal2 542 -914 544 -912 8 s2
rlabel metal1 433 -806 444 -803 1 a2
rlabel metal1 433 -813 444 -810 1 b2
rlabel metal1 466 -808 471 -805 1 p2_inv
rlabel metal1 575 -776 577 -774 1 g2_inv
rlabel metal1 588 -843 593 -841 1 p1_inv
rlabel metal1 652 -730 655 -727 1 temp107
rlabel metal1 590 -837 594 -835 1 p2_inv
rlabel metal1 617 -839 621 -837 1 temp105
rlabel metal1 640 -829 644 -828 1 c1
rlabel metal1 686 -828 688 -826 1 temp106
rlabel metal1 546 -775 552 -772 1 temp108
rlabel metal1 491 -790 493 -788 1 c3
rlabel metal1 520 -812 520 -812 1 gnd
rlabel metal1 530 -731 530 -730 5 vdd
rlabel metal1 559 -804 559 -804 1 gnd
rlabel metal1 568 -731 568 -731 5 vdd
rlabel metal1 595 -766 596 -766 3 vdd
rlabel metal1 677 -756 677 -756 7 gnd
rlabel metal1 660 -858 660 -858 1 gnd
rlabel metal1 651 -785 651 -785 5 vdd
rlabel metal1 605 -860 605 -860 1 gnd
rlabel metal1 595 -779 595 -778 5 vdd
rlabel m2contact 501 -846 501 -846 1 c2
rlabel m2contact 403 -811 409 -808 1 g2_inv
rlabel metal1 658 -772 661 -769 1 g1_inv
rlabel metal1 806 -752 806 -751 5 vdd
rlabel metal1 816 -833 816 -833 1 gnd
rlabel metal1 787 -772 787 -772 5 vdd
rlabel metal1 801 -880 801 -880 3 gnd
rlabel metal1 801 -872 801 -872 3 vdd
rlabel metal2 702 -891 702 -891 1 mid_s3
rlabel metal2 903 -918 905 -916 8 s3
rlabel metal1 861 -853 862 -846 1 c3
rlabel metal1 794 -817 805 -814 1 b3
rlabel metal1 794 -810 805 -807 1 a3
rlabel metal1 765 -816 771 -813 1 g3_inv
rlabel metal1 827 -812 832 -809 1 p3_inv
rlabel metal1 856 -750 856 -749 5 vdd
rlabel metal1 866 -831 866 -831 1 gnd
rlabel metal1 851 -808 855 -806 3 p3_inv
rlabel m2contact 850 -813 852 -812 3 p2_inv
rlabel metal1 880 -810 881 -808 7 temp109
rlabel metal1 898 -755 898 -755 5 vdd
rlabel metal1 907 -828 907 -828 1 gnd
rlabel m2contact 888 -793 891 -790 1 temp101
rlabel metal1 933 -798 935 -796 1 p4
rlabel metal1 1022 -775 1022 -775 5 vdd
rlabel metal1 1031 -848 1031 -848 1 gnd
rlabel metal1 1058 -818 1058 -816 1 temp110
rlabel metal1 993 -836 993 -836 1 gnd
rlabel metal1 1003 -755 1003 -754 5 vdd
rlabel metal1 1010 -818 1010 -818 1 temp109
rlabel metal1 1004 -813 1016 -810 1 temp104
rlabel metal1 964 -814 964 -814 1 temp110
rlabel metal1 1083 -765 1083 -764 5 vdd
rlabel metal1 1093 -846 1093 -846 1 gnd
rlabel metal1 1120 -824 1122 -822 1 temp111
rlabel m2contact 1077 -823 1080 -821 1 g2_inv
rlabel m2contact 1079 -830 1079 -830 1 p3_inv
rlabel metal1 1147 -787 1147 -787 5 vdd
rlabel metal1 1156 -860 1156 -860 1 gnd
rlabel metal1 1163 -831 1169 -828 7 temp112
rlabel metal1 1054 -866 1055 -866 3 vdd
rlabel metal1 1136 -876 1136 -876 7 gnd
rlabel metal1 1113 -892 1115 -889 1 g4_inv
rlabel m2contact 1138 -832 1140 -829 1 g3_inv
rlabel metal1 946 -876 946 -876 3 vdd
rlabel metal1 1019 -885 1019 -885 7 gnd
rlabel metal1 981 -869 984 -867 5 p4
rlabel metal1 946 -910 946 -910 3 vdd
rlabel metal1 1019 -919 1019 -919 7 gnd
rlabel metal1 989 -904 990 -902 7 temp113
rlabel m2contact 981 -903 984 -900 7 g4_inv
rlabel metal1 987 -932 990 -926 1 c4
rlabel m2contact 990 -869 993 -866 5 c0
<< end >>
