* SPICE3 file created from CompleteCircuit.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.global gnd vdd
.option scale=0.09u

M1000 a_81_n604# g1_inv vdd w_75_n617# CMOSP w=40 l=2
+  ad=320 pd=96 as=16860 ps=8216
M1001 c1 mid_s1 s1 w_n309_n731# CMOSP w=20 l=2
+  ad=260 pd=106 as=140 ps=54
M1002 a_n789_n972# a_n814_n972# vdd w_n895_n978# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 p4 a_376_n627# vdd w_326_n648# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 a_832_n935# a_808_n935# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=11150 ps=5990
M1005 b0 a_n779_n520# vdd w_n885_n526# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1006 gnd p1_inv a_n310_n572# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1007 a_n789_n1250# a_n814_n1250# vdd w_n895_n1256# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1008 temp111 a_566_n685# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1009 temp109 p2_inv gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1010 a3 a_n791_n1154# gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1011 a_n883_n1062# b2_in vdd w_n896_n1068# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1012 a_289_n644# b3 vdd w_242_n650# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1013 a_n810_n730# a_n828_n724# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1014 a_n854_n698# a_n878_n730# vdd w_n891_n704# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1015 a_n872_n520# b0_in vdd w_n885_n526# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1016 a_816_n541# c4 vdd w_803_n547# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1017 a_n881_n817# clk a_n881_n785# w_n894_n791# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1018 p3_inv b3 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1019 vdd mid_s0 a_n577_n723# w_n561_n730# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1020 mid_s1 b1 a1 w_n465_n731# CMOSP w=20 l=2
+  ad=240 pd=104 as=200 ps=100
M1021 a_n884_n1186# clk a_n884_n1154# w_n897_n1160# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1022 s0_out a_901_n903# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1023 a1 a_n788_n785# gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1024 a_n814_n1282# a_n832_n1276# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1025 a_129_n695# temp105 gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1026 temp113 c0 vdd w_425_n776# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1027 s1 c1 mid_s1 w_n309_n731# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 p0_inv a0 a_n573_n632# w_n620_n638# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1029 a_882_n628# clk a_882_n660# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1030 c4_out a_909_n541# vdd w_803_n547# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1031 a_876_n903# a_858_n929# vdd w_795_n909# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1032 p0_inv b0 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1033 b3 a3 mid_s3 w_184_n737# CMOSP w=20 l=2
+  ad=200 pd=100 as=240 ps=104
M1034 vdd temp109 a_466_n647# w_434_n655# CMOSP w=40 l=2
+  ad=0 pd=0 as=320 ps=96
M1035 a_n394_n676# b1 g1_inv Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=100 ps=50
M1036 gnd a0 a_n607_n670# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1037 a_814_n628# s3 vdd w_801_n634# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1038 gnd b3 a_195_n761# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1039 b3 a_n789_n1250# vdd w_n895_n1256# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 a_878_n720# a_860_n746# vdd w_797_n726# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1041 a_909_n573# a_884_n541# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1042 a_901_n903# a_876_n903# vdd w_795_n909# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1043 gnd temp109 a_446_n674# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1044 a0 a_n785_n698# vdd w_n891_n704# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1045 vdd b3 a_195_n761# w_224_n742# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1046 a_500_n685# temp104 gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1047 s3_out a_907_n628# vdd w_801_n634# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1048 a2 a_n789_n972# gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1049 p4 a_376_n627# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1050 a_n785_n698# a_n810_n698# vdd w_n891_n704# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1051 a_n850_n639# a_n874_n639# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1052 a_469_n763# temp113 c4 Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=100 ps=50
M1053 s2 c2 a_n76_n731# Gnd CMOSN w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1054 a_n791_n1154# a_n816_n1154# vdd w_n897_n1160# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1055 vdd temp112 a_540_n724# w_534_n737# CMOSP w=40 l=2
+  ad=0 pd=0 as=320 ps=96
M1056 s0_inv s0_out vdd w_949_n910# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1057 a_n781_n607# clk a_n781_n639# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1058 a_907_n660# a_882_n628# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1059 vdd c1 a_129_n657# w_116_n663# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1060 a_78_n671# p1_inv vdd w_65_n677# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1061 a_n858_n1282# clk a_n858_n1250# w_n895_n1256# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1062 a_n806_n607# clk a_n806_n639# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1063 gnd p2_inv temp105 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1064 c4_inv c4_out vdd w_954_n548# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1065 vdd a0 g0_inv w_n620_n638# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1066 a_909_n541# clk a_909_n573# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1067 a_n460_n672# temp100 gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1068 gnd b1 a_n454_n755# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1069 a_n804_n520# a_n822_n546# vdd w_n885_n526# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1070 a_840_n573# a_816_n573# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1071 temp107 a_81_n594# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1072 temp107 a_81_n594# vdd w_75_n617# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1073 a_n856_n914# clk a_n856_n882# w_n893_n888# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1074 a3 a_n791_n1154# vdd w_n897_n1160# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1075 a_n781_n639# a_n806_n607# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 a_n857_n817# a_n881_n817# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1077 a_808_n903# s0 vdd w_795_n909# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1078 a_907_n628# clk a_907_n660# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1079 a_n607_n670# b0 g0_inv Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1080 temp111 a_566_n685# vdd w_553_n663# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1081 a_838_n660# a_814_n660# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1082 a_n858_n1250# a_n882_n1282# vdd w_n895_n1256# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 a_n815_n1062# a_n833_n1088# vdd w_n896_n1068# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1084 a_n859_n1062# a_n883_n1094# vdd w_n896_n1068# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1085 s2_inv s2_out vdd w_950_n727# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1086 a_810_n720# s2 vdd w_797_n726# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1087 a_625_n697# temp111 gnd Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1088 a_903_n720# a_878_n720# vdd w_797_n726# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1089 a_500_n647# temp109 a_500_n685# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1090 a_n878_n730# a0_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1091 s0_out a_901_n903# vdd w_795_n909# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1092 a_n858_n972# a_n882_n1004# vdd w_n895_n978# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1093 temp104 g1_inv a_n205_n609# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=160 ps=56
M1094 s0_inv s0_out gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1095 a_n298_n663# c0 a_n321_n657# Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=100 ps=50
M1096 vdd g1_inv temp104 w_n218_n577# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1097 a_n860_n1186# clk a_n860_n1154# w_n897_n1160# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1098 s2_out a_903_n720# vdd w_797_n726# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1099 a_n810_n698# a_n828_n724# vdd w_n891_n704# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1100 vdd g4_inv c4 w_425_n776# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1101 a_n162_n591# temp102 vdd w_n218_n577# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1102 temp103 a_n310_n572# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1103 c4_inv c4_out gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1104 a_n816_n1154# clk a_n816_n1186# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1105 a_n884_n1186# a3_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1106 s1_out a_900_n806# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1107 a_n788_n817# a_n813_n785# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1108 a_n880_n914# clk a_n880_n882# w_n893_n888# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1109 a_n106_n678# b2 g2_inv Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=100 ps=50
M1110 g0_inv b0 vdd w_n620_n638# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 a_n881_n817# a1_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1112 a_832_n903# a_808_n935# vdd w_795_n909# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1113 a2 a_n789_n972# vdd w_n895_n978# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1114 gnd b2 a_n166_n757# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1115 temp108 g2_inv vdd w_n38_n631# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1116 c0 a_n781_n607# gnd Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1117 a_376_n627# temp109 a_376_n665# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=160 ps=56
M1118 a_n310_n572# p1_inv a_n282_n572# w_n290_n557# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1119 vdd g3_inv temp112 w_612_n665# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1120 a_n828_n724# a_n854_n730# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1121 temp106 a_129_n657# vdd w_116_n663# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1122 a_834_n720# a_810_n752# vdd w_797_n726# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1123 a_n822_n546# a_n848_n552# vdd w_n885_n526# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1124 a_831_n838# clk a_831_n806# w_794_n812# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1125 a_469_n729# c0 temp113 Gnd CMOSN w=20 l=2
+  ad=160 pd=56 as=100 ps=50
M1126 a_901_n903# clk a_901_n935# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1127 a_n882_n972# a2_in vdd w_n895_n978# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1128 a_81_n594# p2_inv a_81_n604# w_75_n617# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1129 a_875_n838# a_857_n832# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1130 a_n779_n520# clk a_n779_n552# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1131 s2_inv s2_out gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1132 a_900_n838# a_875_n806# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1133 a_n813_n785# clk a_n813_n817# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1134 a_n874_n639# clk a_n874_n607# w_n887_n613# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1135 gnd mid_s0 a_n577_n723# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1136 vdd mid_s1 a_n364_n729# w_n348_n736# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1137 a_n831_n811# a_n857_n817# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1138 a_n804_n520# clk a_n804_n552# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1139 a_n667_n749# a0 mid_s0 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=70 ps=34
M1140 a_n205_n609# temp103 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 a_n360_n638# b1 vdd w_n407_n644# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1142 a_909_n541# a_884_n541# vdd w_803_n547# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1143 temp104 temp103 vdd w_n218_n577# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 p1_inv b1 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1145 gnd a0 p0_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 s3_inv s3_out gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1147 gnd a1 a_n394_n676# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1148 a_n790_n1062# clk a_n790_n1094# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1149 a_875_n806# clk a_875_n838# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1150 a_466_n647# temp104 a_446_n674# w_434_n655# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1151 a_n850_n607# a_n874_n639# vdd w_n887_n613# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1152 s2 c2 mid_s2 w_n21_n733# CMOSP w=20 l=2
+  ad=140 pd=54 as=240 ps=104
M1153 a_446_n674# temp104 gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 a_n779_n552# a_n804_n520# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 a_907_n628# a_882_n628# vdd w_801_n634# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1156 a_n857_n785# a_n881_n817# vdd w_n894_n791# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1157 a_n813_n817# a_n831_n811# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 vdd b0 a_n667_n749# w_n638_n730# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1159 a_n832_n998# a_n858_n1004# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1160 temp106 a_129_n657# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1161 a_n789_n972# clk a_n789_n1004# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1162 a_n833_n1088# a_n859_n1094# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1163 mid_s0 a_n667_n749# a0 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1164 a_n856_n914# a_n880_n914# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1165 a_129_n657# temp105 vdd w_116_n663# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 a_n878_n698# a0_in vdd w_n891_n704# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1167 a_n787_n882# clk a_n787_n914# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1168 a_840_n541# a_816_n573# vdd w_803_n547# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1169 a_n814_n972# a_n832_n998# vdd w_n895_n978# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1170 a_n882_n1250# b3_in vdd w_n895_n1256# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1171 a_807_n838# s1 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1172 a_857_n832# a_831_n838# vdd w_794_n812# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1173 vdd p4 temp113 w_425_n776# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 a_n848_n552# clk a_n848_n520# w_n885_n526# CMOSP w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1175 temp105 p1_inv gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 g1_inv b1 vdd w_n407_n644# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1177 a_n816_n1186# a_n834_n1180# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 a1 a_n788_n785# vdd w_n894_n791# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 c1 g0_inv a_n460_n672# Gnd CMOSN w=20 l=2
+  ad=150 pd=80 as=0 ps=0
M1180 a_n860_n1186# a_n884_n1186# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1181 a_n781_n607# a_n806_n607# vdd w_n887_n613# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1182 vdd mid_s2 a_n76_n731# w_n60_n738# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1183 a_500_n647# temp104 vdd w_434_n655# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1184 c0 a_n577_n723# s0 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1185 a_838_n628# a_814_n660# vdd w_801_n634# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1186 vdd b2 a_n166_n757# w_n137_n738# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1187 a_n788_n785# a_n813_n785# vdd w_n894_n791# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1188 a_n72_n640# b2 vdd w_n119_n646# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1189 a_816_n573# clk a_816_n541# w_803_n547# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1190 a_n881_n785# a1_in vdd w_n894_n791# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 c0_inv c0 vdd w_n546_n618# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1192 p2_inv b2 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1193 a_n789_n1250# clk a_n789_n1282# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1194 gnd g4_inv a_469_n763# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 a_n787_n914# a_n812_n882# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 a_n880_n914# b1_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1197 gnd a2 a_n106_n678# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 a_n874_n639# c0_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1199 gnd a3 a_255_n682# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1200 a_814_n660# clk a_814_n628# w_801_n634# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1201 c1 temp100 vdd w_n546_n618# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1202 gnd temp101 a_n298_n663# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 a_n832_n1276# a_n858_n1282# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1204 gnd a_446_n674# temp110 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1205 a_n884_n1154# a3_in vdd w_n897_n1160# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 s3 c3 a_285_n735# Gnd CMOSN w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1207 s0 c0 a_n577_n723# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 a_n162_n619# temp104 a_n162_n591# w_n218_n577# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1209 mid_s3 a_195_n761# a3 Gnd CMOSN w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1210 a_n812_n882# clk a_n812_n914# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1211 s3_inv s3_out vdd w_951_n635# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1212 a_n790_n1094# a_n815_n1062# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 a_n509_n632# p0_inv vdd w_n546_n618# CMOSP w=40 l=2
+  ad=320 pd=96 as=0 ps=0
M1214 a_n832_n998# a_n858_n1004# vdd w_n895_n978# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1215 a_n247_n639# p1_inv temp101 w_n260_n645# CMOSP w=40 l=2
+  ad=320 pd=96 as=200 ps=90
M1216 a_n824_n633# a_n850_n639# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1217 b1 a_n787_n882# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1218 a_875_n806# a_857_n832# vdd w_794_n812# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1219 a_376_n665# temp101 gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 a_n833_n1088# a_n859_n1094# vdd w_n896_n1068# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1221 a_864_n654# a_838_n660# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1222 temp112 temp111 vdd w_612_n665# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 temp101 p1_inv gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1224 vdd temp109 a_500_n647# w_434_n655# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 a_n789_n1004# a_n814_n972# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 a_n321_n657# c0 vdd w_n333_n637# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1227 c0_inv c0 gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1228 a_900_n806# a_875_n806# vdd w_794_n812# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1229 c3 a_285_n735# s3 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1230 a_n813_n785# a_n831_n811# vdd w_n894_n791# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1231 g4_inv temp110 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1232 a_n814_n1250# a_n832_n1276# vdd w_n895_n1256# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1233 a_n162_n619# temp102 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1234 a_n848_n552# a_n872_n552# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1235 a_n856_n882# a_n880_n914# vdd w_n893_n888# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 a_n812_n914# a_n830_n908# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 gnd mid_s1 a_n364_n729# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1238 a_n806_n639# a_n824_n633# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 a_808_n935# clk a_808_n903# w_795_n909# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1240 g2_inv b2 vdd w_n119_n646# CMOSP w=20 l=2
+  ad=160 pd=56 as=0 ps=0
M1241 temp109 p3_inv a_339_n642# w_326_n648# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1242 a_810_n752# clk a_810_n720# w_797_n726# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1243 vdd temp109 a_376_n627# w_326_n648# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1244 p1_inv a1 a_n360_n638# w_n407_n644# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1245 gnd a1 p1_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 vdd a_n27_n650# c3 w_n38_n631# CMOSP w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1247 b1 a_n787_n882# vdd w_n893_n888# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1248 a_n789_n1282# a_n814_n1250# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 gnd p4 a_469_n729# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 a_n828_n724# a_n854_n730# vdd w_n891_n704# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1251 a_n787_n882# a_n812_n882# vdd w_n893_n888# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1252 a_807_n806# s1 vdd w_794_n812# CMOSP w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1253 a_n872_n552# b0_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1254 a_n880_n882# b1_in vdd w_n893_n888# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 a_n858_n1004# clk a_n858_n972# w_n895_n978# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1256 a_860_n746# a_834_n752# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1257 a_n166_n757# a2 mid_s2 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1258 vdd a_446_n674# temp110 w_434_n655# CMOSP w=20 l=2
+  ad=0 pd=0 as=200 ps=100
M1259 a_n816_n1154# a_n834_n1180# vdd w_n897_n1160# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1260 a_n860_n1154# a_n884_n1186# vdd w_n897_n1160# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 s1_out a_900_n806# vdd w_794_n812# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1262 a_834_n752# clk a_834_n720# w_797_n726# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1263 b2 a_n790_n1062# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1264 a_n831_n811# a_n857_n817# vdd w_n894_n791# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1265 c0 a_n781_n607# vdd w_n887_n613# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1266 vdd a1 g1_inv w_n407_n644# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 gnd mid_s2 a_n76_n731# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 temp110 a_500_n647# vdd w_434_n655# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 a_878_n752# a_860_n746# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1270 s1_inv s1_out vdd w_951_n813# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1271 vdd mid_s3 a_285_n735# w_301_n742# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1272 a_n883_n1094# clk a_n883_n1062# w_n896_n1068# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1273 a_n874_n607# c0_in vdd w_n887_n613# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 b0 a_n779_n520# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1275 p2_inv a2 a_n72_n640# w_n119_n646# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1276 a_n858_n1004# a_n882_n1004# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1277 temp103 a_n310_n572# vdd w_n290_n557# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1278 mid_s2 a_n166_n757# a2 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 gnd a_n27_n650# c3 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1280 gnd a2 p2_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 temp100 a_n509_n660# vdd w_n546_n618# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1282 a_255_n682# b3 g3_inv Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1283 s3 c3 mid_s3 w_340_n737# CMOSP w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1284 a_900_n806# clk a_900_n838# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1285 mid_s3 b3 a3 w_184_n737# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1286 a_566_n685# g2_inv a_566_n657# w_553_n663# CMOSP w=40 l=2
+  ad=200 pd=90 as=320 ps=96
M1287 vdd g0_inv c1 w_n546_n618# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1288 a_878_n720# clk a_878_n752# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1289 a_831_n838# a_807_n838# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1290 gnd g2_inv a_566_n685# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1291 a_n854_n730# clk a_n854_n698# w_n891_n704# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1292 a_n872_n552# clk a_n872_n520# w_n885_n526# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1293 a_n804_n552# a_n822_n546# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1294 a_81_n594# g1_inv gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1295 a_n812_n882# a_n830_n908# vdd w_n893_n888# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1296 a_n790_n1062# a_n815_n1062# vdd w_n896_n1068# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1297 a_866_n567# a_840_n573# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1298 gnd temp107 a_36_n641# Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1299 gnd mid_s3 a_285_n735# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 b3 a_n789_n1250# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1301 temp110 a_500_n647# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1302 a_n310_n572# g0_inv gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 a_n830_n908# a_n856_n914# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1304 s1_inv s1_out gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1305 a_n509_n660# c0_inv a_n509_n632# w_n546_n618# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1306 vdd a2 g2_inv w_n119_n646# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 vdd p0_inv a_n247_n639# w_n260_n645# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 a_840_n573# clk a_840_n541# w_803_n547# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1309 a_n858_n1282# a_n882_n1282# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1310 c3 mid_s3 s3 w_340_n737# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 vdd a3 g3_inv w_242_n650# CMOSP w=20 l=2
+  ad=0 pd=0 as=160 ps=56
M1312 vdd a_n321_n657# temp102 w_n333_n637# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1313 s3_out a_907_n628# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1314 a_n509_n660# p0_inv gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1315 a_884_n573# a_866_n567# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1316 a_810_n752# s2 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1317 gnd p0_inv temp101 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1318 a_n857_n817# clk a_n857_n785# w_n894_n791# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1319 a_903_n752# a_878_n720# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1320 c2 a_n76_n731# s2 Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1321 c2 a_n162_n619# vdd w_n218_n577# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1322 a_n791_n1154# clk a_n791_n1186# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1323 a_n806_n607# a_n824_n633# vdd w_n887_n613# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1324 vdd temp101 a_n321_n657# w_n333_n637# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1325 temp100 a_n509_n660# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1326 b2 a_n790_n1062# vdd w_n896_n1068# CMOSP w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1327 b0 a0 mid_s0 w_n678_n725# CMOSP w=20 l=2
+  ad=0 pd=0 as=240 ps=104
M1328 a_838_n660# clk a_838_n628# w_801_n634# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1329 a_n878_n730# clk a_n878_n698# w_n891_n704# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1330 a_882_n660# a_864_n654# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 a0 a_n785_n698# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1332 gnd temp104 a_n162_n619# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 a_n834_n1180# a_n860_n1186# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1334 a_n454_n755# a1 mid_s1 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1335 a_339_n642# p2_inv vdd w_326_n648# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 gnd p3_inv temp109 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1337 a_884_n541# clk a_884_n573# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1338 a_376_n627# temp101 vdd w_326_n648# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 a_903_n720# clk a_903_n752# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1340 a_n779_n520# a_n804_n520# vdd w_n885_n526# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1341 a_n859_n1094# clk a_n859_n1062# w_n896_n1068# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1342 c1 a_n364_n729# s1 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1343 a_834_n752# a_810_n752# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1344 p3_inv a3 a_289_n644# w_242_n650# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1345 a_540_n724# temp110 g4_inv w_534_n737# CMOSP w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1346 a_n830_n908# a_n856_n914# vdd w_n893_n888# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1347 gnd a3 p3_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 mid_s0 b0 a0 w_n678_n725# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1349 a_n815_n1062# clk a_n815_n1094# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1350 b2 a2 mid_s2 w_n177_n733# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 gnd a_n321_n657# temp102 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1352 a_n883_n1094# b2_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1353 a_129_n657# c1 a_129_n695# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1354 a_858_n929# a_832_n935# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1355 a_n832_n1276# a_n858_n1282# vdd w_n895_n1256# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1356 gnd temp112 g4_inv Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 a_n573_n632# b0 vdd w_n620_n638# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 a_816_n573# c4 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1359 s2_out a_903_n720# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1360 vdd b1 a_n454_n755# w_n425_n736# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1361 a_866_n567# a_840_n573# vdd w_803_n547# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1362 a_n882_n1004# a2_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1363 a_n814_n972# clk a_n814_n1004# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1364 mid_s1 a_n454_n755# a1 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1365 a_832_n935# clk a_832_n903# w_795_n909# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1366 s1 c1 a_n364_n729# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 a_876_n935# a_858_n929# gnd Gnd CMOSN w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1368 c0 mid_s0 s0 w_n522_n725# CMOSP w=20 l=2
+  ad=0 pd=0 as=140 ps=54
M1369 a_n824_n633# a_n850_n639# vdd w_n887_n613# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1370 a_195_n761# a3 mid_s3 Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1371 a_814_n660# s3 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1372 mid_s2 b2 a2 w_n177_n733# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1373 a_864_n654# a_838_n660# vdd w_801_n634# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1374 a_901_n935# a_876_n903# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 a_n854_n730# a_n878_n730# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1376 c2 a_n162_n619# gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 a_n785_n698# clk a_n785_n730# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=140 ps=54
M1378 a_n822_n546# a_n848_n552# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1379 temp105 p2_inv a_78_n671# w_65_n677# CMOSP w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1380 a_n7_n623# temp108 a_n27_n650# w_n38_n631# CMOSP w=40 l=2
+  ad=320 pd=96 as=200 ps=90
M1381 a_n791_n1186# a_n816_n1154# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 a_n27_n650# temp108 gnd Gnd CMOSN w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1383 gnd b0 a_n667_n749# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 a_n834_n1180# a_n860_n1186# vdd w_n897_n1160# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1385 a_831_n806# a_807_n838# vdd w_794_n812# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1386 a_876_n903# clk a_876_n935# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1387 a_n882_n1004# clk a_n882_n972# w_n895_n978# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1388 a_n882_n1282# b3_in gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1389 a_n814_n1250# clk a_n814_n1282# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1390 c4 temp113 vdd w_425_n776# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 s0 c0 mid_s0 w_n522_n725# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1392 vdd temp106 a_n7_n623# w_n38_n631# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1393 a_566_n657# p3_inv vdd w_553_n663# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 gnd temp106 a_n27_n650# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 a_n788_n785# clk a_n788_n817# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1396 a_566_n685# p3_inv gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1397 c4_out a_909_n541# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1398 a_n282_n572# g0_inv vdd w_n290_n557# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 a_n785_n730# a_n810_n698# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 a_807_n838# clk a_807_n806# w_794_n812# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1401 a_36_n641# g2_inv temp108 Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1402 temp112 g3_inv a_625_n697# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1403 a_884_n541# a_866_n567# vdd w_803_n547# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1404 gnd p2_inv a_81_n594# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1405 c2 mid_s2 s2 w_n21_n733# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 a_808_n935# s0 gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1407 a_858_n929# a_832_n935# vdd w_795_n909# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1408 a_n815_n1094# a_n833_n1088# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 g3_inv b3 vdd w_242_n650# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1410 a_n850_n639# clk a_n850_n607# w_n887_n613# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1411 a_n859_n1094# a_n883_n1094# gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1412 gnd c0_inv a_n509_n660# Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1413 a_n882_n1282# clk a_n882_n1250# w_n895_n1256# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1414 a_860_n746# a_834_n752# vdd w_797_n726# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1415 a_882_n628# a_864_n654# vdd w_801_n634# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1416 a_n848_n520# a_n872_n552# vdd w_n885_n526# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1417 a_n814_n1004# a_n832_n998# gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1418 a_n810_n698# clk a_n810_n730# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1419 a_857_n832# a_831_n838# gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1420 b1 a1 mid_s1 w_n465_n731# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1421 vdd temp107 temp108 w_n38_n631# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_n810_n698# gnd 0.05fF
C1 c0_inv c0 0.04fF
C2 p1_inv temp101 0.37fF
C3 temp102 a_n321_n657# 0.04fF
C4 w_n21_n733# s2 0.17fF
C5 w_n897_n1160# a_n860_n1186# 0.09fF
C6 w_534_n737# temp112 0.06fF
C7 p0_inv a_n460_n672# 0.00fF
C8 w_n348_n736# mid_s1 0.07fF
C9 w_n895_n978# a2 0.02fF
C10 g0_inv vdd 0.73fF
C11 a_857_n832# gnd 0.05fF
C12 w_434_n655# a_446_n674# 0.09fF
C13 c0_inv gnd 0.03fF
C14 c1 a_n364_n729# 0.10fF
C15 a_n310_n572# g1_inv 0.07fF
C16 w_340_n737# c0 0.01fF
C17 w_797_n726# vdd 0.14fF
C18 temp107 temp106 0.00fF
C19 p3_inv temp110 0.13fF
C20 a3 a_n791_n1154# 0.05fF
C21 w_n897_n1160# a3 0.02fF
C22 g1_inv gnd 0.09fF
C23 a_878_n720# clk 0.03fF
C24 g2_inv a2 0.32fF
C25 p3_inv a_500_n685# 0.01fF
C26 mid_s2 c2 0.27fF
C27 a_858_n929# gnd 0.05fF
C28 temp109 a_376_n627# 0.10fF
C29 a_n810_n698# clk 0.03fF
C30 b1_in a_n880_n914# 0.03fF
C31 w_797_n726# a_878_n720# 0.11fF
C32 c1 b2 0.02fF
C33 w_425_n776# c4 0.04fF
C34 w_n887_n613# a_n781_n607# 0.12fF
C35 b2 a_n790_n1062# 0.05fF
C36 a_814_n660# a_838_n660# 0.03fF
C37 w_949_n910# vdd 0.02fF
C38 w_534_n737# g4_inv 0.02fF
C39 p3_inv vdd 0.05fF
C40 a_857_n832# clk 0.03fF
C41 mid_s0 a_n577_n723# 0.06fF
C42 a_n874_n639# gnd 0.02fF
C43 g0_inv c0_inv 0.12fF
C44 w_242_n650# a3 0.44fF
C45 w_n119_n646# a2 0.44fF
C46 b3 s2 0.08fF
C47 b0 a_n607_n670# 0.01fF
C48 w_794_n812# a_807_n838# 0.09fF
C49 g1_inv g0_inv 0.05fF
C50 a_907_n628# s3_out 0.05fF
C51 b3 a_195_n761# 0.11fF
C52 a_n830_n908# gnd 0.05fF
C53 a_858_n929# clk 0.03fF
C54 w_n333_n637# temp101 0.07fF
C55 a2_in a_n882_n1004# 0.03fF
C56 w_n290_n557# temp103 0.09fF
C57 temp106 vdd 0.24fF
C58 w_n309_n731# s1 0.17fF
C59 w_794_n812# s1_out 0.02fF
C60 g2_inv a_129_n657# 0.01fF
C61 a_n364_n729# c0 0.02fF
C62 w_n38_n631# g2_inv 0.45fF
C63 c4_out c4_inv 0.04fF
C64 a1 vdd 0.12fF
C65 w_n893_n888# a_n880_n914# 0.09fF
C66 w_n885_n526# a_n822_n546# 0.09fF
C67 c2 a_n76_n731# 0.10fF
C68 mid_s2 s2 0.00fF
C69 a_n832_n998# gnd 0.05fF
C70 w_n891_n704# a_n878_n730# 0.09fF
C71 c1 temp105 0.25fF
C72 a_n162_n619# gnd 0.04fF
C73 w_n177_n733# b2 0.10fF
C74 a_n874_n639# clk 0.14fF
C75 s3 mid_s3 0.00fF
C76 a_n364_n729# gnd 0.02fF
C77 w_n546_n618# c1 0.04fF
C78 g1_inv a_n7_n623# 0.01fF
C79 b2 c0 0.04fF
C80 a_n856_n914# a_n830_n908# 0.05fF
C81 w_794_n812# clk 0.14fF
C82 a_n830_n908# clk 0.03fF
C83 c1 c0 0.30fF
C84 w_n620_n638# vdd 0.12fF
C85 w_795_n909# a_876_n903# 0.11fF
C86 w_n895_n1256# vdd 0.14fF
C87 w_116_n663# c1 0.07fF
C88 b2 gnd 0.18fF
C89 w_801_n634# s3 0.07fF
C90 g0_inv a_n509_n632# 0.01fF
C91 a_n832_n998# clk 0.03fF
C92 w_553_n663# a_566_n685# 0.09fF
C93 p0_inv temp100 0.00fF
C94 g1_inv temp106 0.00fF
C95 temp101 vdd 0.16fF
C96 c1 gnd 0.36fF
C97 w_803_n547# c4 0.07fF
C98 mid_s3 vdd 0.12fF
C99 w_612_n665# temp112 0.04fF
C100 a_n858_n1004# a_n832_n998# 0.05fF
C101 w_n60_n738# mid_s2 0.07fF
C102 w_n260_n645# temp102 0.01fF
C103 g1_inv a1 0.32fF
C104 b0 p0_inv 0.02fF
C105 s3_out gnd 0.02fF
C106 w_n887_n613# c0_in 0.07fF
C107 w_116_n663# temp105 0.07fF
C108 w_n546_n618# c0 0.07fF
C109 b0 a_n667_n749# 0.06fF
C110 w_801_n634# vdd 0.14fF
C111 p2_inv b3 0.01fF
C112 temp105 gnd 0.02fF
C113 a_n828_n724# gnd 0.05fF
C114 g0_inv c1 0.10fF
C115 c4 g4_inv 0.54fF
C116 w_n897_n1160# a_n884_n1186# 0.09fF
C117 s0 s1 7.10fF
C118 p0_inv a_n321_n657# 0.01fF
C119 a_81_n594# p2_inv 0.17fF
C120 b0_in gnd 0.02fF
C121 a0 c0 0.17fF
C122 c0 gnd 0.82fF
C123 g1_inv temp101 0.06fF
C124 a_866_n567# gnd 0.05fF
C125 w_n60_n738# a_n76_n731# 0.02fF
C126 w_n407_n644# a1 0.44fF
C127 w_116_n663# gnd 0.01fF
C128 a1_in gnd 0.02fF
C129 b3 s1 0.06fF
C130 a_n310_n572# gnd 0.04fF
C131 g2_inv a_36_n641# 0.01fF
C132 w_340_n737# mid_s3 0.10fF
C133 w_n678_n725# a0 0.24fF
C134 a1 a_n788_n785# 0.05fF
C135 a_807_n838# gnd 0.02fF
C136 a_n828_n724# clk 0.03fF
C137 w_326_n648# p4 0.02fF
C138 g3_inv gnd 0.94fF
C139 temp107 a_81_n594# 0.04fF
C140 w_425_n776# vdd 0.13fF
C141 w_n887_n613# a_n806_n607# 0.11fF
C142 s1_out gnd 0.02fF
C143 w_n546_n618# g0_inv 0.56fF
C144 a_834_n752# clk 0.06fF
C145 a_446_n674# gnd 0.04fF
C146 b0_in clk 0.07fF
C147 a_808_n935# gnd 0.02fF
C148 temp104 temp109 0.47fF
C149 g0_inv c0 0.07fF
C150 w_954_n548# c4_inv 0.02fF
C151 a0_in a_n878_n730# 0.03fF
C152 w_797_n726# a_834_n752# 0.09fF
C153 w_n425_n736# b1 0.15fF
C154 a_866_n567# clk 0.03fF
C155 s0_out gnd 0.02fF
C156 c1 temp106 0.00fF
C157 b1 a2 3.44fF
C158 a1_in clk 0.07fF
C159 w_n218_n577# c2 0.02fF
C160 a2 a_n789_n972# 0.05fF
C161 c3 a_129_n657# 0.01fF
C162 a_n310_n572# g0_inv 0.02fF
C163 g1_inv a_n282_n572# 0.03fF
C164 temp102 p1_inv 0.06fF
C165 w_242_n650# p2_inv 0.32fF
C166 b2_in gnd 0.02fF
C167 w_n38_n631# c3 0.02fF
C168 s3 a_814_n660# 0.03fF
C169 b3 vdd 0.25fF
C170 a1 c1 0.25fF
C171 a_807_n838# clk 0.14fF
C172 g0_inv a0 0.40fF
C173 g0_inv gnd 0.09fF
C174 clk gnd 19.77fF
C175 a_n804_n520# gnd 0.05fF
C176 a_n454_n755# c0 0.22fF
C177 w_950_n727# s2_out 0.07fF
C178 w_n119_n646# g2_inv 0.30fF
C179 temp101 a_n162_n619# 0.00fF
C180 g1_inv a_n205_n609# 0.01fF
C181 w_n885_n526# a_n848_n552# 0.09fF
C182 a_808_n935# clk 0.14fF
C183 a_n813_n785# gnd 0.05fF
C184 a_566_n685# temp111 0.04fF
C185 temp106 temp105 0.01fF
C186 temp110 temp112 0.29fF
C187 w_75_n617# a_81_n594# 0.09fF
C188 mid_s2 vdd 0.12fF
C189 w_n38_n631# temp108 0.13fF
C190 w_n309_n731# c1 0.24fF
C191 a3_in a_n884_n1186# 0.03fF
C192 b2_in clk 0.07fF
C193 a_n856_n914# clk 0.06fF
C194 w_n561_n730# a_n577_n723# 0.02fF
C195 w_n895_n1256# a_n789_n1250# 0.12fF
C196 a_n804_n520# clk 0.03fF
C197 b3_in a_n882_n1282# 0.03fF
C198 w_n897_n1160# vdd 0.14fF
C199 w_n348_n736# vdd 0.11fF
C200 p3_inv gnd 0.95fF
C201 g1_inv a_n27_n650# 0.00fF
C202 p3_inv g3_inv 0.23fF
C203 g0_inv a_n573_n632# 0.01fF
C204 a_n854_n730# a_n828_n724# 0.05fF
C205 w_116_n663# temp106 0.48fF
C206 w_797_n726# clk 0.14fF
C207 a_n858_n1004# clk 0.06fF
C208 p3_inv a_446_n674# 0.05fF
C209 w_803_n547# vdd 0.14fF
C210 a1 c0 0.11fF
C211 w_795_n909# a_832_n935# 0.09fF
C212 a_n813_n785# clk 0.03fF
C213 a_n815_n1062# gnd 0.05fF
C214 w_949_n910# s0_out 0.07fF
C215 temp106 gnd 0.11fF
C216 w_n333_n637# temp102 0.48fF
C217 temp110 g4_inv 0.17fF
C218 a_n814_n1250# gnd 0.05fF
C219 w_n260_n645# p0_inv 0.07fF
C220 w_242_n650# vdd 0.12fF
C221 g1_inv a_81_n594# 0.06fF
C222 w_801_n634# a_907_n628# 0.12fF
C223 p0_inv b1 0.01fF
C224 a0 a1 0.06fF
C225 g2_inv p4 0.01fF
C226 a_864_n654# gnd 0.05fF
C227 w_801_n634# s3_out 0.02fF
C228 w_612_n665# temp111 0.08fF
C229 p1_inv a2 0.67fF
C230 w_803_n547# a_909_n541# 0.12fF
C231 w_n309_n731# c0 0.01fF
C232 b0 mid_s0 0.25fF
C233 w_951_n635# s3_inv 0.02fF
C234 temp109 a_500_n647# 0.10fF
C235 g4_inv vdd 0.02fF
C236 temp103 vdd 0.84fF
C237 a_n860_n1186# a_n834_n1180# 0.05fF
C238 a_n815_n1062# clk 0.03fF
C239 temp101 c0 0.30fF
C240 w_n620_n638# a0 0.44fF
C241 w_553_n663# vdd 0.07fF
C242 w_n465_n731# mid_s1 0.18fF
C243 mid_s3 c0 0.11fF
C244 clk a_n814_n1250# 0.03fF
C245 a_n310_n572# temp101 0.01fF
C246 a_864_n654# clk 0.03fF
C247 temp101 gnd 0.02fF
C248 b2 s0 0.06fF
C249 mid_s3 gnd 0.22fF
C250 temp102 vdd 0.24fF
C251 a_n854_n730# clk 0.06fF
C252 a_285_n735# gnd 0.02fF
C253 a1 a_n454_n755# 0.31fF
C254 a_816_n573# gnd 0.02fF
C255 g2_inv c3 0.06fF
C256 a2 p2_inv 0.17fF
C257 w_n894_n791# vdd 0.14fF
C258 w_n887_n613# a_n824_n633# 0.09fF
C259 w_n620_n638# g0_inv 0.30fF
C260 g2_inv a3 0.34fF
C261 w_n895_n1256# clk 0.14fF
C262 w_434_n655# temp104 0.15fF
C263 w_326_n648# temp109 0.09fF
C264 temp103 g1_inv 0.32fF
C265 w_n465_n731# b1 0.10fF
C266 w_n895_n978# a_n789_n972# 0.12fF
C267 g0_inv temp101 0.00fF
C268 a_376_n627# gnd 0.02fF
C269 w_951_n813# vdd 0.02fF
C270 temp108 g2_inv 0.36fF
C271 b3 a_n789_n1250# 0.05fF
C272 a_n880_n914# gnd 0.02fF
C273 w_n348_n736# a_n364_n729# 0.02fF
C274 p1_inv p0_inv 0.42fF
C275 b2 mid_s2 0.25fF
C276 a2 s1 0.06fF
C277 a_n822_n546# gnd 0.05fF
C278 a_816_n573# clk 0.14fF
C279 g1_inv temp104 0.18fF
C280 temp101 a_n162_n591# 0.01fF
C281 w_n885_n526# a_n872_n552# 0.09fF
C282 c3 a_78_n671# 0.01fF
C283 c1 mid_s2 0.01fF
C284 g1_inv temp102 0.09fF
C285 w_425_n776# c0 0.08fF
C286 a_n882_n1004# gnd 0.02fF
C287 w_801_n634# clk 0.14fF
C288 g2_inv a_566_n685# 0.17fF
C289 a_n831_n811# gnd 0.05fF
C290 s0 c0 0.65fF
C291 a_n880_n914# a_n856_n914# 0.03fF
C292 a_500_n647# temp110 0.04fF
C293 temp101 p3_inv 0.00fF
C294 a_n880_n914# clk 0.14fF
C295 w_794_n812# a_875_n806# 0.11fF
C296 w_65_n677# c3 0.01fF
C297 w_326_n648# p2_inv 0.06fF
C298 a_n822_n546# clk 0.03fF
C299 s0 gnd 0.02fF
C300 w_n896_n1068# vdd 0.14fF
C301 w_n895_n1256# a_n814_n1250# 0.11fF
C302 w_n38_n631# temp107 0.07fF
C303 b3 c0 0.12fF
C304 w_n425_n736# vdd 0.11fF
C305 a2 vdd 0.12fF
C306 p1_inv a_n298_n663# 0.01fF
C307 w_n522_n725# mid_s0 0.10fF
C308 a_n27_n650# gnd 0.04fF
C309 a_n882_n1004# clk 0.14fF
C310 s0 a_808_n935# 0.03fF
C311 w_n218_n577# vdd 0.11fF
C312 p2_inv a_289_n644# 0.01fF
C313 a_n831_n811# clk 0.03fF
C314 temp112 a_625_n697# 0.00fF
C315 a_n833_n1088# gnd 0.05fF
C316 b3 gnd 0.05fF
C317 w_n177_n733# mid_s2 0.18fF
C318 a_n882_n1004# a_n858_n1004# 0.03fF
C319 b3 g3_inv 0.32fF
C320 a_n162_n619# temp104 0.17fF
C321 a_n832_n1276# gnd 0.05fF
C322 mid_s2 c0 0.01fF
C323 w_n333_n637# p0_inv 0.01fF
C324 p0_inv a_n509_n660# 0.02fF
C325 temp102 a_n162_n619# 0.02fF
C326 s0 clk 0.07fF
C327 a_81_n594# gnd 0.04fF
C328 w_184_n737# a3 0.24fF
C329 w_224_n742# b3 0.13fF
C330 w_n894_n791# a_n788_n785# 0.12fF
C331 mid_s2 gnd 0.22fF
C332 w_n348_n736# c0 0.02fF
C333 w_434_n655# a_500_n647# 0.11fF
C334 a_n878_n730# gnd 0.02fF
C335 w_n38_n631# vdd 0.11fF
C336 w_n895_n978# a2_in 0.07fF
C337 w_801_n634# a_864_n654# 0.09fF
C338 g2_inv temp109 0.02fF
C339 a_814_n660# gnd 0.02fF
C340 a_n833_n1088# clk 0.03fF
C341 w_803_n547# a_866_n567# 0.09fF
C342 clk a_n832_n1276# 0.03fF
C343 w_954_n548# c4_out 0.07fF
C344 w_n218_n577# g1_inv 0.09fF
C345 s2 a_810_n752# 0.03fF
C346 temp112 gnd 0.15fF
C347 g3_inv temp112 0.11fF
C348 b1 a_n394_n676# 0.01fF
C349 w_n137_n738# a_n166_n757# 0.02fF
C350 w_326_n648# vdd 0.09fF
C351 mid_s3 a_285_n735# 0.06fF
C352 a_n76_n731# c0 0.04fF
C353 a_n878_n730# clk 0.14fF
C354 p0_inv vdd 0.09fF
C355 c3 a3 0.01fF
C356 c4 temp113 0.10fF
C357 a_814_n660# clk 0.14fF
C358 w_n887_n613# a_n850_n639# 0.09fF
C359 c0 g4_inv 0.04fF
C360 a_n76_n731# gnd 0.02fF
C361 b3 p3_inv 0.02fF
C362 w_242_n650# g3_inv 0.04fF
C363 w_n897_n1160# clk 0.14fF
C364 w_n38_n631# g1_inv 0.02fF
C365 b1 mid_s1 0.31fF
C366 a1 s0 0.06fF
C367 temp103 a_n310_n572# 0.04fF
C368 temp106 a_n27_n650# 0.02fF
C369 g2_inv p2_inv 0.11fF
C370 w_301_n742# vdd 0.11fF
C371 w_n895_n978# a_n814_n972# 0.11fF
C372 p1_inv a_n321_n657# 0.01fF
C373 a_n282_n572# temp101 0.00fF
C374 w_803_n547# clk 0.14fF
C375 w_n885_n526# b0 0.02fF
C376 g4_inv gnd 0.09fF
C377 g2_inv a_81_n604# 0.02fF
C378 a2 a_n364_n729# 0.14fF
C379 temp102 c0 0.00fF
C380 w_n218_n577# a_n162_n619# 0.09fF
C381 a_831_n838# a_857_n832# 0.05fF
C382 w_65_n677# p1_inv 0.06fF
C383 a_875_n806# gnd 0.05fF
C384 p0_inv c0_inv 0.25fF
C385 w_n119_n646# p2_inv 0.02fF
C386 temp107 g2_inv 0.32fF
C387 w_950_n727# vdd 0.02fF
C388 a_n509_n660# temp100 0.04fF
C389 g1_inv p0_inv 0.06fF
C390 w_n896_n1068# b2 0.02fF
C391 temp102 gnd 0.11fF
C392 a_n577_n723# c0 0.10fF
C393 w_n894_n791# a1_in 0.07fF
C394 s1_out s1_inv 0.04fF
C395 b2 a2 5.50fF
C396 b1 a_n787_n882# 0.05fF
C397 a_876_n903# gnd 0.05fF
C398 temp104 a_446_n674# 0.17fF
C399 w_797_n726# a_903_n720# 0.12fF
C400 w_n896_n1068# a_n790_n1062# 0.12fF
C401 c1 a2 0.08fF
C402 w_n895_n1256# b3 0.02fF
C403 a_832_n935# a_858_n929# 0.05fF
C404 w_n638_n730# a_n667_n749# 0.02fF
C405 a3_in gnd 0.02fF
C406 a_n848_n552# clk 0.06fF
C407 w_n895_n1256# a_n832_n1276# 0.09fF
C408 a_n577_n723# gnd 0.02fF
C409 w_n895_n978# vdd 0.14fF
C410 a_875_n806# clk 0.03fF
C411 w_n561_n730# mid_s0 0.07fF
C412 w_242_n650# p3_inv 0.02fF
C413 a_n878_n730# a_n854_n730# 0.03fF
C414 b3 mid_s3 0.32fF
C415 a3 s2 0.06fF
C416 w_n887_n613# vdd 0.14fF
C417 b2 a_n166_n757# 0.26fF
C418 a_n857_n817# clk 0.06fF
C419 s0_out s0_inv 0.04fF
C420 w_794_n812# a_831_n838# 0.09fF
C421 w_65_n677# p2_inv 0.37fF
C422 a3 a_195_n761# 0.10fF
C423 a_876_n903# clk 0.03fF
C424 w_n333_n637# a_n321_n657# 0.11fF
C425 g2_inv vdd 0.23fF
C426 w_951_n813# s1_out 0.07fF
C427 w_75_n617# g2_inv 0.01fF
C428 w_n894_n791# clk 0.14fF
C429 w_n407_n644# p0_inv 0.02fF
C430 w_553_n663# p3_inv 0.06fF
C431 c2 s2 0.35fF
C432 c1 a_129_n657# 0.10fF
C433 a3_in clk 0.07fF
C434 c0_in a_n874_n639# 0.03fF
C435 w_n894_n791# a_n813_n785# 0.11fF
C436 b0 vdd 0.19fF
C437 w_n177_n733# a2 0.24fF
C438 w_n425_n736# c0 0.01fF
C439 a2 c0 0.50fF
C440 p1_inv c3 0.00fF
C441 w_n119_n646# vdd 0.12fF
C442 w_n290_n557# p1_inv 0.07fF
C443 p3_inv temp104 0.01fF
C444 a_n884_n1186# a_n860_n1186# 0.03fF
C445 a_n859_n1094# clk 0.06fF
C446 w_795_n909# a_901_n903# 0.12fF
C447 clk a_n858_n1282# 0.06fF
C448 a_n816_n1154# gnd 0.05fF
C449 a2 gnd 0.14fF
C450 w_949_n910# s0_inv 0.02fF
C451 w_801_n634# a_814_n660# 0.09fF
C452 a_n781_n607# c0 0.05fF
C453 g1_inv g2_inv 0.02fF
C454 p0_inv c1 0.17fF
C455 a_n166_n757# c0 0.04fF
C456 w_803_n547# a_816_n573# 0.09fF
C457 a_500_n647# gnd 0.02fF
C458 p1_inv c2 0.01fF
C459 w_n21_n733# mid_s2 0.10fF
C460 w_n260_n645# p1_inv 0.47fF
C461 p1_inv b1 0.02fF
C462 g3_inv temp111 0.21fF
C463 w_n896_n1068# b2_in 0.07fF
C464 w_n887_n613# a_n874_n639# 0.09fF
C465 w_65_n677# vdd 0.02fF
C466 b3 s0 0.06fF
C467 a_834_n752# a_860_n746# 0.05fF
C468 w_116_n663# a_129_n657# 0.11fF
C469 p2_inv c3 0.14fF
C470 a_n816_n1154# clk 0.03fF
C471 w_n894_n791# a1 0.02fF
C472 w_n896_n1068# clk 0.14fF
C473 w_951_n635# vdd 0.02fF
C474 b0_in a_n872_n552# 0.03fF
C475 w_n638_n730# b0 0.07fF
C476 temp103 temp101 0.01fF
C477 a_n850_n639# a_n824_n633# 0.05fF
C478 p2_inv a3 0.01fF
C479 a1 a_n577_n723# 0.60fF
C480 a_129_n657# gnd 0.06fF
C481 mid_s0 vdd 0.12fF
C482 w_n895_n978# a_n832_n998# 0.09fF
C483 w_n893_n888# a_n787_n882# 0.12fF
C484 w_n891_n704# a_n785_n698# 0.12fF
C485 p4 vdd 0.13fF
C486 mid_s1 s1 0.00fF
C487 w_n546_n618# p0_inv 0.06fF
C488 w_n425_n736# a_n454_n755# 0.02fF
C489 a_860_n746# gnd 0.05fF
C490 a_909_n541# c4_out 0.05fF
C491 temp101 temp104 0.01fF
C492 w_n893_n888# b1 0.02fF
C493 a_n872_n552# gnd 0.02fF
C494 w_534_n737# temp110 0.06fF
C495 a1_in a_n881_n817# 0.03fF
C496 temp102 temp101 0.07fF
C497 p0_inv c0 0.28fF
C498 a_884_n541# gnd 0.05fF
C499 c3 s3 0.35fF
C500 a3 s1 0.06fF
C501 a_n881_n817# gnd 0.02fF
C502 a_807_n838# a_831_n838# 0.03fF
C503 a_n779_n520# b0 0.05fF
C504 a0 p0_inv 0.17fF
C505 p0_inv gnd 0.61fF
C506 w_534_n737# vdd 0.02fF
C507 w_n896_n1068# a_n815_n1062# 0.11fF
C508 p3_inv a_500_n647# 0.05fF
C509 a_860_n746# clk 0.03fF
C510 a0 a_n667_n749# 0.14fF
C511 a_n872_n552# clk 0.14fF
C512 mid_s1 vdd 0.12fF
C513 g2_inv b2 0.27fF
C514 w_n895_n1256# a_n858_n1282# 0.09fF
C515 a_n848_n552# a_n822_n546# 0.05fF
C516 g2_inv a_376_n665# 0.01fF
C517 a_884_n541# clk 0.03fF
C518 w_797_n726# a_860_n746# 0.09fF
C519 c1 g2_inv 0.00fF
C520 c3 vdd 0.07fF
C521 w_n290_n557# vdd 0.09fF
C522 a_n881_n817# clk 0.14fF
C523 a_808_n935# a_832_n935# 0.03fF
C524 w_425_n776# g4_inv 0.10fF
C525 a_n883_n1094# gnd 0.02fF
C526 w_795_n909# vdd 0.14fF
C527 a3 vdd 0.12fF
C528 a_831_n838# clk 0.06fF
C529 c0_in gnd 0.02fF
C530 g0_inv p0_inv 0.05fF
C531 w_242_n650# b3 0.14fF
C532 a_n882_n1282# gnd 0.02fF
C533 w_n119_n646# b2 0.14fF
C534 a_n857_n817# a_n831_n811# 0.05fF
C535 temp102 a_n205_n609# 0.01fF
C536 w_n897_n1160# a_n791_n1154# 0.12fF
C537 a_832_n935# clk 0.06fF
C538 g2_inv temp105 0.00fF
C539 w_n894_n791# a_n831_n811# 0.09fF
C540 temp106 a_129_n657# 0.04fF
C541 w_n38_n631# temp106 0.06fF
C542 b2_in a_n883_n1094# 0.03fF
C543 w_n260_n645# vdd 0.02fF
C544 b1 vdd 0.22fF
C545 w_n893_n888# b1_in 0.07fF
C546 w_326_n648# p3_inv 0.06fF
C547 s3_out s3_inv 0.04fF
C548 mid_s2 a_n76_n731# 0.06fF
C549 w_n891_n704# a0_in 0.07fF
C550 s1 s2 6.42fF
C551 a_n883_n1094# clk 0.14fF
C552 w_n887_n613# c0 0.02fF
C553 p2_inv temp109 0.02fF
C554 a_n834_n1180# gnd 0.05fF
C555 s3 s2 5.40fF
C556 clk a_n882_n1282# 0.14fF
C557 c0_in clk 0.07fF
C558 w_n218_n577# temp101 0.03fF
C559 w_n546_n618# temp100 0.09fF
C560 p1_inv p2_inv 0.28fF
C561 w_n290_n557# g1_inv 0.01fF
C562 w_116_n663# g2_inv 0.02fF
C563 c4 s3 3.18fF
C564 w_954_n548# vdd 0.02fF
C565 w_795_n909# a_858_n929# 0.09fF
C566 w_340_n737# c3 0.24fF
C567 g2_inv gnd 0.09fF
C568 b0 c0 0.02fF
C569 g2_inv g3_inv 0.00fF
C570 a_n806_n607# gnd 0.05fF
C571 g3_inv a_255_n682# 0.01fF
C572 w_n891_n704# vdd 0.14fF
C573 g1_inv temp108 0.01fF
C574 p0_inv a1 0.05fF
C575 temp112 g4_inv 0.02fF
C576 a_882_n628# gnd 0.05fF
C577 g1_inv c2 0.05fF
C578 a_n834_n1180# clk 0.03fF
C579 w_n895_n978# clk 0.14fF
C580 w_951_n635# s3_out 0.07fF
C581 w_n678_n725# b0 0.10fF
C582 g1_inv b1 0.26fF
C583 a1 a_n667_n749# 0.66fF
C584 b0 a0 0.91fF
C585 b0 gnd 0.05fF
C586 a_n859_n1094# a_n833_n1088# 0.05fF
C587 w_n895_n978# a_n858_n1004# 0.09fF
C588 w_n887_n613# clk 0.14fF
C589 w_n893_n888# a_n812_n882# 0.11fF
C590 a_810_n752# a_834_n752# 0.03fF
C591 w_65_n677# temp105 0.05fF
C592 w_n891_n704# a_n810_n698# 0.11fF
C593 mid_s1 a_n364_n729# 0.06fF
C594 w_612_n665# vdd 0.05fF
C595 w_n620_n638# p0_inv 0.02fF
C596 a_n321_n657# c0 0.10fF
C597 a_n806_n607# clk 0.03fF
C598 a_n858_n1282# a_n832_n1276# 0.05fF
C599 w_326_n648# temp101 0.43fF
C600 temp113 c0 0.11fF
C601 g0_inv temp100 0.31fF
C602 w_950_n727# s2_inv 0.02fF
C603 a_882_n628# clk 0.03fF
C604 a_840_n573# a_866_n567# 0.05fF
C605 w_n897_n1160# a3_in 0.07fF
C606 p0_inv temp101 0.08fF
C607 a_n321_n657# gnd 0.06fF
C608 p1_inv vdd 0.63fF
C609 a_810_n752# gnd 0.02fF
C610 a2 s0 0.06fF
C611 b0 g0_inv 0.26fF
C612 w_n60_n738# vdd 0.11fF
C613 c1 mid_s1 0.27fF
C614 mid_s0 c0 0.42fF
C615 w_n896_n1068# a_n833_n1088# 0.09fF
C616 w_n407_n644# b1 0.14fF
C617 s2_out gnd 0.02fF
C618 a_n162_n619# c2 0.04fF
C619 c4_out gnd 0.02fF
C620 p4 c0 0.30fF
C621 b2 a3 10.24fF
C622 temp106 a_36_n641# 0.01fF
C623 g2_inv p3_inv 0.28fF
C624 w_301_n742# mid_s3 0.07fF
C625 w_n895_n1256# a_n882_n1282# 0.09fF
C626 c1 c3 0.00fF
C627 w_n561_n730# vdd 0.11fF
C628 w_326_n648# a_376_n627# 0.11fF
C629 w_434_n655# temp109 0.14fF
C630 w_n678_n725# mid_s0 0.18fF
C631 temp103 temp102 0.00fF
C632 w_301_n742# a_285_n735# 0.02fF
C633 w_184_n737# c0 0.01fF
C634 mid_s0 gnd 0.22fF
C635 w_n465_n731# a1 0.24fF
C636 a0 mid_s0 0.40fF
C637 w_n885_n526# vdd 0.14fF
C638 a_810_n752# clk 0.14fF
C639 w_n893_n888# vdd 0.14fF
C640 p4 gnd 0.16fF
C641 temp106 g2_inv 0.16fF
C642 g3_inv p4 0.07fF
C643 a2 mid_s2 0.40fF
C644 w_797_n726# a_810_n752# 0.09fF
C645 a_840_n573# clk 0.06fF
C646 temp102 temp104 0.24fF
C647 p2_inv vdd 0.84fF
C648 temp102 a_n247_n639# 0.01fF
C649 c3 temp105 0.05fF
C650 c1 c2 0.03fF
C651 g1_inv p1_inv 0.05fF
C652 w_n38_n631# a_n27_n650# 0.09fF
C653 w_75_n617# p2_inv 0.07fF
C654 w_n897_n1160# a_n816_n1154# 0.11fF
C655 b1 c1 0.20fF
C656 b3_in gnd 0.02fF
C657 b2 a_n106_n678# 0.01fF
C658 mid_s1 c0 0.05fF
C659 w_797_n726# s2_out 0.02fF
C660 w_n894_n791# a_n857_n817# 0.09fF
C661 w_n522_n725# c0 0.24fF
C662 w_n333_n637# vdd 0.07fF
C663 c3 c0 0.05fF
C664 temp107 vdd 0.84fF
C665 w_794_n812# a_900_n806# 0.12fF
C666 temp106 a_78_n671# 0.01fF
C667 w_116_n663# c3 0.01fF
C668 mid_s1 gnd 0.22fF
C669 a3 c0 0.05fF
C670 w_75_n617# temp107 0.09fF
C671 w_n290_n557# a_n310_n572# 0.09fF
C672 w_951_n813# s1_inv 0.02fF
C673 temp111 temp112 0.00fF
C674 s3 vdd 0.08fF
C675 temp101 g2_inv 0.00fF
C676 c3 gnd 0.12fF
C677 w_n620_n638# b0 0.14fF
C678 c3 g3_inv 0.01fF
C679 temp110 vdd 0.04fF
C680 b3_in clk 0.07fF
C681 a3 gnd 0.03fF
C682 g1_inv p2_inv 0.29fF
C683 w_n407_n644# p1_inv 0.02fF
C684 a_n824_n633# gnd 0.05fF
C685 a3 g3_inv 0.35fF
C686 c2 c0 0.50fF
C687 w_65_n677# temp106 0.01fF
C688 s2_out s2_inv 0.04fF
C689 b1 c0 0.14fF
C690 w_795_n909# a_808_n935# 0.09fF
C691 p3_inv p4 0.05fF
C692 c0_inv a_n509_n660# 0.17fF
C693 a_n860_n1186# clk 0.06fF
C694 w_795_n909# s0_out 0.02fF
C695 w_n218_n577# temp103 0.07fF
C696 a_n874_n639# a_n850_n639# 0.03fF
C697 w_n290_n557# g0_inv 0.06fF
C698 w_n895_n978# a_n882_n1004# 0.09fF
C699 w_801_n634# a_882_n628# 0.11fF
C700 w_75_n617# vdd 0.09fF
C701 w_434_n655# temp110 0.05fF
C702 w_n893_n888# a_n830_n908# 0.09fF
C703 b1 gnd 0.05fF
C704 g1_inv temp107 0.04fF
C705 g2_inv a_376_n627# 0.01fF
C706 w_n885_n526# a_n779_n520# 0.12fF
C707 w_n891_n704# a_n828_n724# 0.09fF
C708 w_795_n909# clk 0.14fF
C709 w_553_n663# temp111 0.02fF
C710 p1_inv b2 0.19fF
C711 w_803_n547# a_884_n541# 0.11fF
C712 a_566_n685# gnd 0.04fF
C713 a_n824_n633# clk 0.03fF
C714 w_n218_n577# temp104 0.13fF
C715 a_n106_n678# gnd 0.01fF
C716 w_n218_n577# temp102 0.06fF
C717 p1_inv c1 0.00fF
C718 w_340_n737# s3 0.17fF
C719 w_434_n655# vdd 0.16fF
C720 p0_inv a_n360_n638# 0.01fF
C721 s2 c0 0.05fF
C722 w_n137_n738# vdd 0.11fF
C723 c4 c0 0.03fF
C724 a_838_n660# clk 0.06fF
C725 a_816_n573# a_840_n573# 0.03fF
C726 w_794_n812# s1 0.07fF
C727 w_n891_n704# a0 0.02fF
C728 w_n896_n1068# a_n859_n1094# 0.09fF
C729 a3 p3_inv 0.17fF
C730 s2 gnd 0.02fF
C731 g1_inv vdd 0.35fF
C732 w_n638_n730# vdd 0.11fF
C733 p1_inv temp105 0.02fF
C734 a_n872_n552# a_n848_n552# 0.03fF
C735 w_75_n617# g1_inv 0.11fF
C736 b1 a_n454_n755# 0.10fF
C737 a1 mid_s1 0.40fF
C738 temp106 c3 0.05fF
C739 g2_inv a_n27_n650# 0.07fF
C740 c4 gnd 0.26fF
C741 b2 p2_inv 0.02fF
C742 g2_inv b3 0.00fF
C743 w_n895_n1256# b3_in 0.07fF
C744 c1 p2_inv 0.00fF
C745 w_184_n737# mid_s3 0.18fF
C746 b3 a_255_n682# 0.01fF
C747 p1_inv c0 0.06fF
C748 w_612_n665# g3_inv 0.07fF
C749 w_n60_n738# c0 0.01fF
C750 w_224_n742# a_195_n761# 0.02fF
C751 a_n881_n817# a_n857_n817# 0.03fF
C752 a0 a_n785_n698# 0.05fF
C753 w_n891_n704# clk 0.14fF
C754 s2 clk 0.07fF
C755 a_n310_n572# p1_inv 0.17fF
C756 a_900_n806# s1_out 0.05fF
C757 temp109 gnd 0.04fF
C758 w_794_n812# vdd 0.14fF
C759 temp108 temp106 0.24fF
C760 w_n897_n1160# a_n834_n1180# 0.09fF
C761 p3_inv a_566_n685# 0.02fF
C762 b1_in gnd 0.02fF
C763 p0_inv a_n247_n639# 0.01fF
C764 w_n309_n731# mid_s1 0.10fF
C765 b2 s1 0.06fF
C766 temp102 p0_inv 0.06fF
C767 p1_inv gnd 0.79fF
C768 w_n894_n791# a_n881_n817# 0.09fF
C769 c4 clk 0.07fF
C770 w_797_n726# s2 0.07fF
C771 a_376_n627# p4 0.04fF
C772 temp109 a_446_n674# 0.02fF
C773 w_n407_n644# vdd 0.12fF
C774 w_n885_n526# b0_in 0.07fF
C775 c1 s1 0.35fF
C776 p2_inv temp105 0.17fF
C777 w_425_n776# temp113 0.11fF
C778 a2_in gnd 0.02fF
C779 b1 a1 4.08fF
C780 a_n884_n1186# gnd 0.02fF
C781 a_838_n660# a_864_n654# 0.05fF
C782 w_n290_n557# temp101 0.02fF
C783 c3 mid_s3 0.28fF
C784 a_901_n903# s0_out 0.05fF
C785 a3 mid_s3 0.40fF
C786 c3 a_285_n735# 0.10fF
C787 a2 a_n166_n757# 0.10fF
C788 b1_in clk 0.07fF
C789 p1_inv g0_inv 0.27fF
C790 w_794_n812# a_857_n832# 0.09fF
C791 w_n546_n618# a_n509_n660# 0.09fF
C792 mid_s0 s0 0.00fF
C793 w_425_n776# p4 0.07fF
C794 b2 vdd 0.19fF
C795 w_242_n650# g2_inv 0.01fF
C796 w_n333_n637# c0 0.07fF
C797 a2_in clk 0.07fF
C798 p2_inv gnd 0.21fF
C799 c1 vdd 0.12fF
C800 p2_inv g3_inv 0.00fF
C801 a_n884_n1186# clk 0.14fF
C802 w_n260_n645# temp101 0.05fF
C803 c0 a_469_n763# 0.02fF
C804 a_n812_n882# gnd 0.05fF
C805 w_n407_n644# g1_inv 0.04fF
C806 s1 c0 0.05fF
C807 a_n883_n1094# a_n859_n1094# 0.03fF
C808 g1_inv a_n162_n619# 0.04fF
C809 w_n333_n637# gnd 0.01fF
C810 a_n509_n660# gnd 0.04fF
C811 w_n893_n888# a_n856_n914# 0.09fF
C812 w_n885_n526# clk 0.14fF
C813 p3_inv temp109 0.18fF
C814 w_n885_n526# a_n804_n520# 0.11fF
C815 s3 c0 0.01fF
C816 w_n891_n704# a_n854_n730# 0.09fF
C817 w_553_n663# g2_inv 0.10fF
C818 a_n814_n972# gnd 0.05fF
C819 w_n893_n888# clk 0.14fF
C820 w_184_n737# b3 0.10fF
C821 s1 a_807_n838# 0.03fF
C822 a_n882_n1282# a_n858_n1282# 0.03fF
C823 a_n850_n639# clk 0.06fF
C824 w_n137_n738# b2 0.20fF
C825 s1 gnd 0.02fF
C826 a0_in gnd 0.02fF
C827 w_801_n634# a_838_n660# 0.09fF
C828 s3 gnd 0.02fF
C829 w_n546_n618# vdd 0.14fF
C830 a_n812_n882# clk 0.03fF
C831 p1_inv temp106 0.00fF
C832 w_803_n547# a_840_n573# 0.09fF
C833 w_n522_n725# s0 0.17fF
C834 temp110 gnd 0.26fF
C835 g3_inv temp110 0.37fF
C836 w_n21_n733# c2 0.24fF
C837 w_803_n547# c4_out 0.02fF
C838 g0_inv a_n509_n660# 0.05fF
C839 p1_inv a1 0.17fF
C840 c0 vdd 0.63fF
C841 a_n814_n972# clk 0.03fF
C842 a_446_n674# temp110 0.04fF
C843 w_n896_n1068# a_n883_n1094# 0.09fF
C844 w_116_n663# vdd 0.07fF
C845 w_795_n909# s0 0.07fF
C846 a3 s0 0.06fF
C847 a_n27_n650# c3 0.04fF
C848 s1 clk 0.07fF
C849 a0_in clk 0.07fF
C850 a0 vdd 0.12fF
C851 vdd gnd 2.08fF
C852 c3 b3 0.02fF
C853 p2_inv p3_inv 0.38fF
C854 c4 a_816_n573# 0.03fF
C855 s3 clk 0.07fF
C856 g3_inv vdd 0.57fF
C857 a_903_n720# s2_out 0.05fF
C858 temp113 g4_inv 0.33fF
C859 b3 a3 8.83fF
C860 w_n546_n618# c0_inv 0.12fF
C861 a_878_n720# gnd 0.05fF
C862 temp101 temp109 0.24fF
C863 b1 s0 0.06fF
C864 temp106 p2_inv 0.06fF
C865 g2_inv a_n72_n640# 0.01fF
C866 temp108 a_n27_n650# 0.17fF
C867 w_n137_n738# c0 0.01fF
C868 w_224_n742# vdd 0.11fF
C869 gnd Gnd 10.30fF
C870 vdd Gnd 10.21fF
C871 a_n789_n1250# Gnd 0.17fF
C872 a_n814_n1250# Gnd 0.15fF
C873 a_n832_n1276# Gnd 0.17fF
C874 a_n858_n1282# Gnd 0.19fF
C875 a_n882_n1282# Gnd 0.05fF
C876 clk Gnd 7.58fF
C877 b3_in Gnd 0.13fF
C878 a_n791_n1154# Gnd 0.17fF
C879 a_n816_n1154# Gnd 0.15fF
C880 a_n834_n1180# Gnd 0.17fF
C881 a_n860_n1186# Gnd 0.19fF
C882 a_n884_n1186# Gnd 0.05fF
C883 a3_in Gnd 0.13fF
C884 a_n790_n1062# Gnd 0.17fF
C885 a_n815_n1062# Gnd 0.15fF
C886 a_n833_n1088# Gnd 0.17fF
C887 a_n859_n1094# Gnd 0.19fF
C888 a_n883_n1094# Gnd 0.16fF
C889 b2_in Gnd 0.10fF
C890 a_n789_n972# Gnd 0.17fF
C891 a_n814_n972# Gnd 0.15fF
C892 a_n832_n998# Gnd 0.17fF
C893 a_n858_n1004# Gnd 0.19fF
C894 a_n882_n1004# Gnd 0.16fF
C895 a2_in Gnd 0.10fF
C896 s0_inv Gnd 0.02fF
C897 s0_out Gnd 0.22fF
C898 a_901_n903# Gnd 0.17fF
C899 a_876_n903# Gnd 0.15fF
C900 a_858_n929# Gnd 0.17fF
C901 a_832_n935# Gnd 0.19fF
C902 a_808_n935# Gnd 0.16fF
C903 a_n787_n882# Gnd 0.17fF
C904 a_n812_n882# Gnd 0.15fF
C905 a_n830_n908# Gnd 0.17fF
C906 a_n856_n914# Gnd 0.19fF
C907 a_n880_n914# Gnd 0.16fF
C908 b1_in Gnd 0.13fF
C909 s1_inv Gnd 0.02fF
C910 s1_out Gnd 0.23fF
C911 a_900_n806# Gnd 0.17fF
C912 a_875_n806# Gnd 0.15fF
C913 a_857_n832# Gnd 0.17fF
C914 a_831_n838# Gnd 0.19fF
C915 a_807_n838# Gnd 0.16fF
C916 s2_inv Gnd 0.02fF
C917 a_n788_n785# Gnd 0.17fF
C918 a_n813_n785# Gnd 0.15fF
C919 a_n831_n811# Gnd 0.17fF
C920 a_n857_n817# Gnd 0.19fF
C921 a_n881_n817# Gnd 0.16fF
C922 a1_in Gnd 0.13fF
C923 s2_out Gnd 0.21fF
C924 g4_inv Gnd 0.55fF
C925 c0 Gnd 3.10fF
C926 temp113 Gnd 0.24fF
C927 a_285_n735# Gnd 0.38fF
C928 a_195_n761# Gnd 0.38fF
C929 a_903_n720# Gnd 0.17fF
C930 a_878_n720# Gnd 0.15fF
C931 a_860_n746# Gnd 0.17fF
C932 a_834_n752# Gnd 0.19fF
C933 a_810_n752# Gnd 0.16fF
C934 mid_s3 Gnd 1.09fF
C935 s2 Gnd 5.55fF
C936 a_n76_n731# Gnd 0.38fF
C937 a_n166_n757# Gnd 0.38fF
C938 s3_inv Gnd 0.03fF
C939 temp112 Gnd 0.04fF
C940 temp111 Gnd 0.03fF
C941 s3_out Gnd 0.21fF
C942 a_566_n685# Gnd 0.18fF
C943 temp110 Gnd 0.28fF
C944 a_500_n647# Gnd 0.18fF
C945 a_907_n628# Gnd 0.17fF
C946 a_882_n628# Gnd 0.15fF
C947 a_864_n654# Gnd 0.17fF
C948 a_838_n660# Gnd 0.19fF
C949 a_814_n660# Gnd 0.05fF
C950 s3 Gnd 0.45fF
C951 c2 Gnd 0.75fF
C952 mid_s2 Gnd 1.09fF
C953 s1 Gnd 8.75fF
C954 a_n364_n729# Gnd 0.38fF
C955 a_n454_n755# Gnd 0.38fF
C956 mid_s1 Gnd 1.09fF
C957 s0 Gnd 11.79fF
C958 a_n577_n723# Gnd 0.38fF
C959 a_n667_n749# Gnd 0.28fF
C960 a_446_n674# Gnd 0.18fF
C961 p4 Gnd 0.54fF
C962 a_376_n627# Gnd 0.00fF
C963 temp109 Gnd 0.41fF
C964 temp104 Gnd 0.59fF
C965 g3_inv Gnd 2.47fF
C966 mid_s0 Gnd 0.22fF
C967 a_129_n657# Gnd 0.12fF
C968 temp105 Gnd 0.31fF
C969 p3_inv Gnd 0.02fF
C970 a3 Gnd 5.85fF
C971 b3 Gnd 6.17fF
C972 c4_inv Gnd 0.03fF
C973 c3 Gnd 0.24fF
C974 a_n27_n650# Gnd 0.18fF
C975 p2_inv Gnd 0.70fF
C976 a_n785_n698# Gnd 0.17fF
C977 a_n810_n698# Gnd 0.15fF
C978 a_n828_n724# Gnd 0.17fF
C979 a_n854_n730# Gnd 0.19fF
C980 a_n878_n730# Gnd 0.03fF
C981 a0_in Gnd 0.10fF
C982 a2 Gnd 4.25fF
C983 b2 Gnd 4.54fF
C984 g2_inv Gnd 2.53fF
C985 temp106 Gnd 0.95fF
C986 temp108 Gnd 0.14fF
C987 a_81_n594# Gnd 0.18fF
C988 temp107 Gnd 0.20fF
C989 a_n162_n619# Gnd 0.17fF
C990 a_n321_n657# Gnd 0.18fF
C991 temp101 Gnd 1.45fF
C992 c1 Gnd 0.48fF
C993 temp100 Gnd 0.19fF
C994 a1 Gnd 3.17fF
C995 b1 Gnd 3.41fF
C996 a_n509_n660# Gnd 0.02fF
C997 c0_inv Gnd 0.11fF
C998 p0_inv Gnd 0.78fF
C999 a0 Gnd 2.47fF
C1000 a_n781_n607# Gnd 0.17fF
C1001 a_n806_n607# Gnd 0.15fF
C1002 a_n824_n633# Gnd 0.17fF
C1003 a_n850_n639# Gnd 0.19fF
C1004 a_n874_n639# Gnd 0.03fF
C1005 c0_in Gnd 0.09fF
C1006 g0_inv Gnd 0.57fF
C1007 p1_inv Gnd 0.48fF
C1008 temp102 Gnd 0.29fF
C1009 g1_inv Gnd 1.56fF
C1010 a_n310_n572# Gnd 0.01fF
C1011 c4_out Gnd 0.21fF
C1012 temp103 Gnd 0.49fF
C1013 a_909_n541# Gnd 0.17fF
C1014 a_884_n541# Gnd 0.15fF
C1015 a_866_n567# Gnd 0.17fF
C1016 a_840_n573# Gnd 0.19fF
C1017 a_816_n573# Gnd 0.05fF
C1018 c4 Gnd 0.06fF
C1019 b0 Gnd 1.99fF
C1020 a_n779_n520# Gnd 0.17fF
C1021 a_n804_n520# Gnd 0.15fF
C1022 a_n822_n546# Gnd 0.17fF
C1023 a_n848_n552# Gnd 0.19fF
C1024 a_n872_n552# Gnd 0.04fF
C1025 b0_in Gnd 0.12fF
C1026 w_n895_n1256# Gnd 0.80fF
C1027 w_n897_n1160# Gnd 0.84fF
C1028 w_n896_n1068# Gnd 0.84fF
C1029 w_n895_n978# Gnd 0.87fF
C1030 w_949_n910# Gnd 0.80fF
C1031 w_795_n909# Gnd 4.56fF
C1032 w_n893_n888# Gnd 0.77fF
C1033 w_951_n813# Gnd 0.80fF
C1034 w_794_n812# Gnd 4.56fF
C1035 w_950_n727# Gnd 0.80fF
C1036 w_797_n726# Gnd 0.05fF
C1037 w_534_n737# Gnd 1.78fF
C1038 w_425_n776# Gnd 2.12fF
C1039 w_n894_n791# Gnd 0.90fF
C1040 w_340_n737# Gnd 1.06fF
C1041 w_301_n742# Gnd 0.84fF
C1042 w_224_n742# Gnd 0.84fF
C1043 w_184_n737# Gnd 1.06fF
C1044 w_n21_n733# Gnd 1.06fF
C1045 w_n60_n738# Gnd 0.84fF
C1046 w_n137_n738# Gnd 0.84fF
C1047 w_n177_n733# Gnd 1.06fF
C1048 w_n309_n731# Gnd 1.06fF
C1049 w_n348_n736# Gnd 0.84fF
C1050 w_n425_n736# Gnd 0.84fF
C1051 w_n465_n731# Gnd 1.06fF
C1052 w_n522_n725# Gnd 1.06fF
C1053 w_n561_n730# Gnd 0.84fF
C1054 w_n638_n730# Gnd 0.16fF
C1055 w_n678_n725# Gnd 0.13fF
C1056 w_951_n635# Gnd 0.58fF
C1057 w_801_n634# Gnd 4.56fF
C1058 w_612_n665# Gnd 1.09fF
C1059 w_553_n663# Gnd 2.17fF
C1060 w_434_n655# Gnd 2.78fF
C1061 w_326_n648# Gnd 2.44fF
C1062 w_116_n663# Gnd 1.82fF
C1063 w_65_n677# Gnd 1.72fF
C1064 w_n891_n704# Gnd 4.56fF
C1065 w_242_n650# Gnd 1.98fF
C1066 w_75_n617# Gnd 0.16fF
C1067 w_n38_n631# Gnd 0.65fF
C1068 w_n119_n646# Gnd 0.71fF
C1069 w_n260_n645# Gnd 1.64fF
C1070 w_n333_n637# Gnd 0.89fF
C1071 w_n407_n644# Gnd 0.19fF
C1072 w_n546_n618# Gnd 4.13fF
C1073 w_n620_n638# Gnd 0.71fF
C1074 w_954_n548# Gnd 0.58fF
C1075 w_803_n547# Gnd 4.56fF
C1076 w_n218_n577# Gnd 0.39fF
C1077 w_n887_n613# Gnd 4.56fF
C1078 w_n290_n557# Gnd 2.17fF
C1079 w_n885_n526# Gnd 4.56fF


Vdd vdd gnd 'SUPPLY'

vclk clk gnd pulse 0 1.8 0ns 10ps 10ps 10ns 20ns

* INPUTS HERE
Va0 a0_in gnd 1.8
Va1 a1_in gnd 0
Va3 a2_in gnd 1.8
Va4 a3_in gnd 0

Vb0 b0_in gnd 1.8
Vb1 b1_in gnd 1.8
Vb2 b2_in gnd 1.8
Vb3 b3_in gnd 0

Vc0 c0_in gnd 0

.ic v(a0)=0
.ic v(a1)=0
.ic v(c0)=0
.ic v(a2)=0
.ic v(a3)=0
.ic v(b0)=0
.ic v(b1)=0
.ic v(b2)=0
.ic v(b3)=0
.ic v(a0_in)=0
.ic v(a1_in)=0
.ic v(a2_in)=0
.ic v(a3_in)=0
.ic v(b0_in)=0
.ic v(b1_in)=0
.ic v(b2_in)=0
.ic v(b3_in)=0
.ic v(s0)=0
* .ic v(s0_out)=0
.ic v(s1)=0
* .ic v(s1_out)=0
.ic v(s2)=0
* .ic v(s2_out)=0
.ic v(s3)=0
* .ic v(s3_out)=0
.ic v(c4)=0
* .ic v(c4_out)=0

* tpd from b0 to s3
.measure tran tpd_rise
+ TRIG v(b0) VAL='0.5*SUPPLY' RISE=1 
+ TARG v(s3) VAL='0.5*SUPPLY' RISE=1

.measure tran tpd_fall
+ TRIG v(b0) VAL='0.5*SUPPLY' FALL=1 
+ TARG v(s3) VAL='0.5*SUPPLY' FALL=1

.measure tran tpd param = '(tpd_rise + tpd_fall)/2'

.tran 100p 400ns

.control
set hcopypscolor = 0
set color0=white 
set color1=black 

run

set curplottitle="2023112005_CLA_Adder"

plot v(a0), v(a1)+2, v(a2)+4, v(a3)+6, v(clk)+8
plot v(b0), v(b1)+2, v(b2)+4, v(b3)+6, v(c0)+8, v(clk)+10
plot v(s3_out)+6, v(s2_out)+4, v(s1_out)+2, v(s0_out), v(c4_out)+8, v(clk)+10
.endc