magic
tech scmos
timestamp 1731351952
<< nwell >>
rect -24 64 10 86
rect -24 34 29 64
rect 4 32 29 34
<< ntransistor >>
rect -13 12 -11 22
rect -3 12 -1 22
rect 15 16 17 26
<< ptransistor >>
rect -13 40 -11 80
rect -3 40 -1 80
rect 15 38 17 58
<< ndiffusion >>
rect -18 16 -13 22
rect -14 12 -13 16
rect -11 18 -9 22
rect -5 18 -3 22
rect -11 12 -3 18
rect -1 16 4 22
rect 10 20 15 26
rect 14 16 15 20
rect 17 22 18 26
rect 17 16 22 22
rect -1 12 0 16
<< pdiffusion >>
rect -14 76 -13 80
rect -18 40 -13 76
rect -11 40 -3 80
rect -1 44 4 80
rect -1 40 0 44
rect 14 54 15 58
rect 10 38 15 54
rect 17 42 22 58
rect 17 38 18 42
<< ndcontact >>
rect -18 12 -14 16
rect -9 18 -5 22
rect 10 16 14 20
rect 18 22 22 26
rect 0 12 4 16
<< pdcontact >>
rect -18 76 -14 80
rect 0 40 4 44
rect 10 54 14 58
rect 18 38 22 42
<< polysilicon >>
rect -13 80 -11 83
rect -3 80 -1 83
rect 15 58 17 61
rect -13 22 -11 40
rect -3 22 -1 40
rect 15 26 17 38
rect 15 13 17 16
rect -13 9 -11 12
rect -3 9 -1 12
<< polycontact >>
rect -17 23 -13 27
rect -7 29 -3 33
rect 11 27 15 31
<< metal1 >>
rect -24 87 13 90
rect -18 80 -15 87
rect 10 68 13 87
rect 10 65 29 68
rect 10 58 13 65
rect -24 30 -7 33
rect 1 31 4 40
rect 19 31 22 38
rect 1 28 11 31
rect -24 24 -17 27
rect 1 26 4 28
rect 19 28 29 31
rect 19 26 22 28
rect -8 23 4 26
rect -8 22 -5 23
rect -18 8 -15 12
rect 1 8 4 12
rect 10 8 13 16
rect -24 5 13 8
<< labels >>
rlabel metal1 -17 88 -17 89 5 vdd
rlabel metal1 -7 7 -7 7 1 gnd
rlabel metal1 -23 25 -22 26 3 in1
rlabel metal1 -21 31 -21 31 3 in2
rlabel metal1 21 30 21 30 1 out
<< end >>
