magic
tech scmos
timestamp 1731382820
<< nwell >>
rect -195 75 -82 107
<< ntransistor >>
rect -184 38 -182 58
rect -150 38 -148 58
rect -119 44 -117 64
rect -95 44 -93 64
<< ptransistor >>
rect -184 81 -182 101
rect -174 81 -172 101
rect -150 81 -148 101
rect -140 81 -138 101
rect -119 81 -117 101
rect -95 81 -93 101
<< ndiffusion >>
rect -189 42 -184 58
rect -185 38 -184 42
rect -182 54 -181 58
rect -182 38 -177 54
rect -155 42 -150 58
rect -151 38 -150 42
rect -148 54 -147 58
rect -148 38 -143 54
rect -124 48 -119 64
rect -120 44 -119 48
rect -117 60 -116 64
rect -117 44 -112 60
rect -100 48 -95 64
rect -96 44 -95 48
rect -93 60 -92 64
rect -93 44 -88 60
<< pdiffusion >>
rect -185 97 -184 101
rect -189 81 -184 97
rect -182 81 -174 101
rect -172 85 -167 101
rect -172 81 -171 85
rect -151 97 -150 101
rect -155 81 -150 97
rect -148 81 -140 101
rect -138 85 -133 101
rect -138 81 -137 85
rect -120 97 -119 101
rect -124 81 -119 97
rect -117 85 -112 101
rect -117 81 -116 85
rect -96 97 -95 101
rect -100 81 -95 97
rect -93 85 -88 101
rect -93 81 -92 85
<< ndcontact >>
rect -189 38 -185 42
rect -181 54 -177 58
rect -155 38 -151 42
rect -147 54 -143 58
rect -124 44 -120 48
rect -116 60 -112 64
rect -100 44 -96 48
rect -92 60 -88 64
<< pdcontact >>
rect -189 97 -185 101
rect -171 81 -167 85
rect -155 97 -151 101
rect -137 81 -133 85
rect -124 97 -120 101
rect -116 81 -112 85
rect -100 97 -96 101
rect -92 81 -88 85
<< polysilicon >>
rect -184 101 -182 105
rect -174 101 -172 105
rect -150 101 -148 105
rect -140 101 -138 105
rect -119 101 -117 105
rect -95 101 -93 105
rect -184 58 -182 81
rect -174 62 -172 81
rect -150 58 -148 81
rect -140 62 -138 81
rect -119 64 -117 81
rect -95 64 -93 81
rect -119 41 -117 44
rect -95 41 -93 44
rect -184 35 -182 38
rect -150 35 -148 38
<< polycontact >>
rect -188 70 -184 74
rect -178 63 -174 67
rect -154 70 -150 74
rect -144 63 -140 67
rect -123 68 -119 72
rect -99 68 -95 72
<< metal1 >>
rect -189 108 -97 111
rect -189 101 -186 108
rect -155 101 -152 108
rect -124 101 -121 108
rect -100 101 -97 108
rect -197 70 -188 73
rect -170 73 -167 81
rect -170 70 -154 73
rect -136 72 -133 81
rect -116 72 -112 81
rect -199 63 -178 66
rect -170 58 -167 70
rect -136 69 -123 72
rect -159 63 -144 66
rect -136 58 -133 69
rect -116 68 -99 72
rect -92 71 -88 81
rect -92 68 -82 71
rect -116 64 -112 68
rect -92 64 -88 68
rect -177 55 -167 58
rect -143 55 -133 58
rect -124 39 -121 44
rect -100 39 -97 44
rect -189 35 -186 38
rect -155 35 -152 38
rect -140 36 -97 39
rect -140 35 -137 36
rect -189 32 -137 35
<< labels >>
rlabel metal1 -194 72 -194 72 1 d
rlabel metal1 -198 64 -197 65 3 clk
rlabel metal1 -87 69 -87 69 7 out
rlabel metal1 -116 37 -116 37 1 gnd
rlabel metal1 -162 71 -162 71 1 mid
rlabel metal1 -157 64 -157 64 1 clk
rlabel metal1 -135 66 -135 66 1 q
rlabel metal1 -188 109 -188 109 5 vdd
<< end >>
