magic
tech scmos
timestamp 1731616366
<< nwell >>
rect -314 361 -237 383
rect -197 377 -165 396
rect -332 351 -237 361
rect -219 371 -165 377
rect -332 331 -280 351
rect -219 343 -167 371
rect -332 329 -308 331
rect -500 296 -468 315
rect -500 290 -446 296
rect -498 262 -446 290
rect -428 280 -351 302
rect -229 283 -195 335
rect -178 323 -144 329
rect -178 297 -122 323
rect -147 291 -122 297
rect -428 270 -333 280
rect -521 242 -487 248
rect -543 216 -487 242
rect -543 210 -518 216
rect -470 202 -436 254
rect -385 250 -333 270
rect -357 248 -333 250
rect -104 249 -70 269
rect -104 247 -36 249
rect -123 243 -36 247
rect -123 217 -15 243
rect -123 215 -98 217
rect -39 211 -15 217
rect -4 237 30 259
rect -4 207 49 237
rect -663 161 -605 183
rect -403 174 -342 206
rect 24 205 49 207
rect 55 205 89 237
rect -263 195 -229 200
rect -300 189 -229 195
rect -322 163 -229 189
rect -663 151 -556 161
rect -322 157 -297 163
rect -734 110 -673 142
rect -639 131 -556 151
rect -611 129 -556 131
rect -540 122 -479 154
rect -263 148 -229 163
rect -208 132 -147 164
rect -23 133 29 167
rect -75 92 -7 124
rect -379 57 -318 58
rect -227 57 -166 58
rect -688 54 -627 55
rect -528 54 -467 55
rect -688 43 -590 54
rect -528 43 -430 54
rect -379 46 -281 57
rect -227 46 -129 57
rect -688 23 -556 43
rect -528 23 -396 43
rect -379 26 -247 46
rect -227 26 -95 46
rect -624 11 -556 23
rect -464 11 -396 23
rect -315 14 -247 26
rect -163 14 -95 26
rect -624 2 -590 11
rect -464 2 -430 11
rect -315 5 -281 14
rect -163 5 -129 14
<< ntransistor >>
rect -159 382 -149 384
rect -155 364 -145 366
rect -155 354 -145 356
rect -321 313 -319 323
rect -260 319 -258 339
rect -250 319 -248 339
rect -303 309 -301 319
rect -293 309 -291 319
rect -516 301 -506 303
rect -520 283 -510 285
rect -520 273 -510 275
rect -417 238 -415 258
rect -407 238 -405 258
rect -218 261 -216 271
rect -208 261 -206 271
rect -167 265 -165 285
rect -157 265 -155 285
rect -136 275 -134 285
rect -374 228 -372 238
rect -364 228 -362 238
rect -346 232 -344 242
rect -531 194 -529 204
rect -510 184 -508 204
rect -500 184 -498 204
rect -459 180 -457 190
rect -449 180 -447 190
rect -111 199 -109 209
rect -93 195 -91 205
rect -83 195 -81 205
rect -652 135 -650 145
rect -392 157 -390 167
rect -383 157 -381 167
rect -355 158 -353 168
rect -59 185 -57 205
rect -49 185 -47 205
rect -28 195 -26 205
rect 7 185 9 195
rect 17 185 19 195
rect 35 189 37 199
rect 66 173 68 193
rect 76 173 78 193
rect -628 109 -626 119
rect -618 109 -616 119
rect -600 113 -598 123
rect -310 141 -308 151
rect -289 131 -287 151
rect -279 131 -277 151
rect 41 154 51 156
rect 41 144 51 146
rect -723 93 -721 103
rect -714 93 -712 103
rect -686 94 -684 104
rect -579 97 -577 117
rect -569 97 -567 117
rect -252 126 -250 136
rect -242 126 -240 136
rect -197 116 -195 126
rect -529 105 -527 115
rect -520 105 -518 115
rect -492 106 -490 116
rect -169 115 -167 125
rect -160 115 -158 125
rect -677 62 -675 72
rect -668 62 -666 72
rect -640 61 -638 71
rect -613 66 -611 76
rect -603 66 -601 76
rect -579 55 -577 75
rect -569 55 -567 75
rect -517 62 -515 72
rect -508 62 -506 72
rect -480 61 -478 71
rect -453 66 -451 76
rect -443 66 -441 76
rect -419 55 -417 75
rect -409 55 -407 75
rect -368 65 -366 75
rect -359 65 -357 75
rect -331 64 -329 74
rect -304 69 -302 79
rect -294 69 -292 79
rect -270 58 -268 78
rect -260 58 -258 78
rect -216 65 -214 75
rect -207 65 -205 75
rect -179 64 -177 74
rect -152 69 -150 79
rect -142 69 -140 79
rect -118 58 -116 78
rect -108 58 -106 78
rect -64 60 -62 80
rect -54 60 -52 80
rect -30 60 -28 80
rect -20 60 -18 80
<< ptransistor >>
rect -191 382 -171 384
rect -321 335 -319 355
rect -303 337 -301 377
rect -293 337 -291 377
rect -260 357 -258 377
rect -250 357 -248 377
rect -213 364 -173 366
rect -213 354 -173 356
rect -494 301 -474 303
rect -492 283 -452 285
rect -417 276 -415 296
rect -407 276 -405 296
rect -492 273 -452 275
rect -531 216 -529 236
rect -510 222 -508 242
rect -500 222 -498 242
rect -459 208 -457 248
rect -449 208 -447 248
rect -374 256 -372 296
rect -364 256 -362 296
rect -218 289 -216 329
rect -208 289 -206 329
rect -167 303 -165 323
rect -157 303 -155 323
rect -346 254 -344 274
rect -136 297 -134 317
rect -111 221 -109 241
rect -93 223 -91 263
rect -83 223 -81 263
rect -59 223 -57 243
rect -49 223 -47 243
rect -392 180 -390 200
rect -383 180 -381 200
rect -355 180 -353 200
rect -28 217 -26 237
rect 7 213 9 253
rect 17 213 19 253
rect -652 157 -650 177
rect -723 116 -721 136
rect -714 116 -712 136
rect -686 116 -684 136
rect -628 137 -626 177
rect -618 137 -616 177
rect -600 135 -598 155
rect -579 135 -577 155
rect -569 135 -567 155
rect -310 163 -308 183
rect -289 169 -287 189
rect -279 169 -277 189
rect -252 154 -250 194
rect -242 154 -240 194
rect 35 211 37 231
rect 66 211 68 231
rect 76 211 78 231
rect -529 128 -527 148
rect -520 128 -518 148
rect -492 128 -490 148
rect -197 138 -195 158
rect -169 138 -167 158
rect -160 138 -158 158
rect -17 154 23 156
rect -17 144 23 146
rect -64 98 -62 118
rect -54 98 -52 118
rect -30 98 -28 118
rect -20 98 -18 118
rect -677 29 -675 49
rect -668 29 -666 49
rect -640 29 -638 49
rect -613 8 -611 48
rect -603 8 -601 48
rect -579 17 -577 37
rect -569 17 -567 37
rect -517 29 -515 49
rect -508 29 -506 49
rect -480 29 -478 49
rect -453 8 -451 48
rect -443 8 -441 48
rect -419 17 -417 37
rect -409 17 -407 37
rect -368 32 -366 52
rect -359 32 -357 52
rect -331 32 -329 52
rect -304 11 -302 51
rect -294 11 -292 51
rect -270 20 -268 40
rect -260 20 -258 40
rect -216 32 -214 52
rect -207 32 -205 52
rect -179 32 -177 52
rect -152 11 -150 51
rect -142 11 -140 51
rect -118 20 -116 40
rect -108 20 -106 40
<< ndiffusion >>
rect -155 385 -149 389
rect -159 384 -149 385
rect -159 381 -149 382
rect -159 377 -153 381
rect -155 367 -149 371
rect -155 366 -145 367
rect -155 362 -145 364
rect -151 358 -145 362
rect -155 356 -145 358
rect -155 353 -145 354
rect -155 349 -149 353
rect -322 319 -321 323
rect -326 313 -321 319
rect -319 317 -314 323
rect -261 335 -260 339
rect -265 319 -260 335
rect -258 319 -250 339
rect -248 323 -243 339
rect -248 319 -247 323
rect -319 313 -318 317
rect -308 313 -303 319
rect -304 309 -303 313
rect -301 315 -299 319
rect -295 315 -293 319
rect -301 309 -293 315
rect -291 313 -286 319
rect -291 309 -290 313
rect -516 304 -510 308
rect -516 303 -506 304
rect -516 300 -506 301
rect -512 296 -506 300
rect -516 286 -510 290
rect -520 285 -510 286
rect -520 281 -510 283
rect -520 277 -514 281
rect -520 275 -510 277
rect -520 272 -510 273
rect -516 268 -510 272
rect -422 242 -417 258
rect -418 238 -417 242
rect -415 238 -407 258
rect -405 254 -404 258
rect -405 238 -400 254
rect -223 265 -218 271
rect -219 261 -218 265
rect -216 267 -214 271
rect -210 267 -208 271
rect -216 261 -208 267
rect -206 265 -201 271
rect -172 269 -167 285
rect -168 265 -167 269
rect -165 265 -157 285
rect -155 281 -154 285
rect -155 265 -150 281
rect -141 279 -136 285
rect -137 275 -136 279
rect -134 281 -133 285
rect -134 275 -129 281
rect -206 261 -205 265
rect -379 232 -374 238
rect -375 228 -374 232
rect -372 234 -370 238
rect -366 234 -364 238
rect -372 228 -364 234
rect -362 232 -357 238
rect -351 236 -346 242
rect -347 232 -346 236
rect -344 238 -343 242
rect -344 232 -339 238
rect -362 228 -361 232
rect -532 200 -531 204
rect -536 194 -531 200
rect -529 198 -524 204
rect -529 194 -528 198
rect -511 200 -510 204
rect -515 184 -510 200
rect -508 184 -500 204
rect -498 188 -493 204
rect -112 205 -111 209
rect -498 184 -497 188
rect -464 184 -459 190
rect -460 180 -459 184
rect -457 186 -455 190
rect -451 186 -449 190
rect -457 180 -449 186
rect -447 184 -442 190
rect -447 180 -446 184
rect -116 199 -111 205
rect -109 203 -104 209
rect -109 199 -108 203
rect -98 199 -93 205
rect -94 195 -93 199
rect -91 201 -89 205
rect -85 201 -83 205
rect -91 195 -83 201
rect -81 199 -76 205
rect -81 195 -80 199
rect -657 139 -652 145
rect -653 135 -652 139
rect -650 141 -649 145
rect -650 135 -645 141
rect -393 163 -392 167
rect -397 157 -392 163
rect -390 163 -388 167
rect -384 163 -383 167
rect -390 157 -383 163
rect -381 161 -376 167
rect -381 157 -380 161
rect -360 162 -355 168
rect -356 158 -355 162
rect -353 162 -348 168
rect -353 158 -352 162
rect -64 189 -59 205
rect -60 185 -59 189
rect -57 185 -49 205
rect -47 201 -46 205
rect -47 185 -42 201
rect -33 199 -28 205
rect -29 195 -28 199
rect -26 201 -25 205
rect -26 195 -21 201
rect 2 189 7 195
rect 6 185 7 189
rect 9 191 11 195
rect 15 191 17 195
rect 9 185 17 191
rect 19 189 24 195
rect 30 193 35 199
rect 34 189 35 193
rect 37 195 38 199
rect 37 189 42 195
rect 19 185 20 189
rect 61 177 66 193
rect 65 173 66 177
rect 68 173 76 193
rect 78 189 79 193
rect 78 173 83 189
rect -633 113 -628 119
rect -629 109 -628 113
rect -626 115 -624 119
rect -620 115 -618 119
rect -626 109 -618 115
rect -616 113 -611 119
rect -605 117 -600 123
rect -601 113 -600 117
rect -598 119 -597 123
rect -598 113 -593 119
rect -311 147 -310 151
rect -315 141 -310 147
rect -308 145 -303 151
rect -308 141 -307 145
rect -290 147 -289 151
rect -294 131 -289 147
rect -287 131 -279 151
rect -277 135 -272 151
rect 41 157 47 161
rect 41 156 51 157
rect 41 152 51 154
rect 45 148 51 152
rect 41 146 51 148
rect 41 143 51 144
rect 41 139 47 143
rect -277 131 -276 135
rect -616 109 -615 113
rect -724 99 -723 103
rect -728 93 -723 99
rect -721 99 -719 103
rect -715 99 -714 103
rect -721 93 -714 99
rect -712 97 -707 103
rect -712 93 -711 97
rect -691 98 -686 104
rect -687 94 -686 98
rect -684 98 -679 104
rect -684 94 -683 98
rect -584 101 -579 117
rect -580 97 -579 101
rect -577 97 -569 117
rect -567 113 -566 117
rect -257 130 -252 136
rect -253 126 -252 130
rect -250 132 -248 136
rect -244 132 -242 136
rect -250 126 -242 132
rect -240 130 -235 136
rect -240 126 -239 130
rect -202 120 -197 126
rect -198 116 -197 120
rect -195 120 -190 126
rect -195 116 -194 120
rect -174 119 -169 125
rect -567 97 -562 113
rect -530 111 -529 115
rect -534 105 -529 111
rect -527 111 -525 115
rect -521 111 -520 115
rect -527 105 -520 111
rect -518 109 -513 115
rect -518 105 -517 109
rect -497 110 -492 116
rect -493 106 -492 110
rect -490 110 -485 116
rect -170 115 -169 119
rect -167 121 -166 125
rect -162 121 -160 125
rect -167 115 -160 121
rect -158 121 -157 125
rect -158 115 -153 121
rect -490 106 -489 110
rect -682 66 -677 72
rect -678 62 -677 66
rect -675 66 -668 72
rect -675 62 -673 66
rect -669 62 -668 66
rect -666 68 -665 72
rect -614 72 -613 76
rect -666 62 -661 68
rect -641 67 -640 71
rect -645 61 -640 67
rect -638 67 -637 71
rect -638 61 -633 67
rect -618 66 -613 72
rect -611 70 -603 76
rect -611 66 -609 70
rect -605 66 -603 70
rect -601 72 -600 76
rect -601 66 -596 72
rect -580 71 -579 75
rect -584 55 -579 71
rect -577 55 -569 75
rect -567 59 -562 75
rect -522 66 -517 72
rect -518 62 -517 66
rect -515 66 -508 72
rect -515 62 -513 66
rect -509 62 -508 66
rect -506 68 -505 72
rect -454 72 -453 76
rect -506 62 -501 68
rect -481 67 -480 71
rect -567 55 -566 59
rect -485 61 -480 67
rect -478 67 -477 71
rect -478 61 -473 67
rect -458 66 -453 72
rect -451 70 -443 76
rect -451 66 -449 70
rect -445 66 -443 70
rect -441 72 -440 76
rect -441 66 -436 72
rect -420 71 -419 75
rect -424 55 -419 71
rect -417 55 -409 75
rect -407 59 -402 75
rect -373 69 -368 75
rect -369 65 -368 69
rect -366 69 -359 75
rect -366 65 -364 69
rect -360 65 -359 69
rect -357 71 -356 75
rect -305 75 -304 79
rect -357 65 -352 71
rect -332 70 -331 74
rect -407 55 -406 59
rect -336 64 -331 70
rect -329 70 -328 74
rect -329 64 -324 70
rect -309 69 -304 75
rect -302 73 -294 79
rect -302 69 -300 73
rect -296 69 -294 73
rect -292 75 -291 79
rect -292 69 -287 75
rect -271 74 -270 78
rect -275 58 -270 74
rect -268 58 -260 78
rect -258 62 -253 78
rect -221 69 -216 75
rect -217 65 -216 69
rect -214 69 -207 75
rect -214 65 -212 69
rect -208 65 -207 69
rect -205 71 -204 75
rect -153 75 -152 79
rect -205 65 -200 71
rect -180 70 -179 74
rect -258 58 -257 62
rect -184 64 -179 70
rect -177 70 -176 74
rect -177 64 -172 70
rect -157 69 -152 75
rect -150 73 -142 79
rect -150 69 -148 73
rect -144 69 -142 73
rect -140 75 -139 79
rect -140 69 -135 75
rect -119 74 -118 78
rect -123 58 -118 74
rect -116 58 -108 78
rect -106 62 -101 78
rect -106 58 -105 62
rect -69 64 -64 80
rect -65 60 -64 64
rect -62 60 -54 80
rect -52 76 -51 80
rect -52 60 -47 76
rect -35 64 -30 80
rect -31 60 -30 64
rect -28 60 -20 80
rect -18 76 -17 80
rect -18 60 -13 76
<< pdiffusion >>
rect -191 385 -175 389
rect -191 384 -171 385
rect -191 381 -171 382
rect -187 377 -171 381
rect -326 339 -321 355
rect -322 335 -321 339
rect -319 351 -318 355
rect -319 335 -314 351
rect -308 341 -303 377
rect -304 337 -303 341
rect -301 337 -293 377
rect -291 373 -290 377
rect -291 337 -286 373
rect -261 373 -260 377
rect -265 357 -260 373
rect -258 361 -250 377
rect -258 357 -256 361
rect -252 357 -250 361
rect -248 373 -247 377
rect -248 357 -243 373
rect -213 367 -177 371
rect -213 366 -173 367
rect -213 356 -173 364
rect -213 353 -173 354
rect -209 349 -173 353
rect -219 325 -218 329
rect -490 304 -474 308
rect -494 303 -474 304
rect -494 300 -474 301
rect -494 296 -478 300
rect -418 292 -417 296
rect -488 286 -452 290
rect -492 285 -452 286
rect -492 275 -452 283
rect -422 276 -417 292
rect -415 280 -407 296
rect -415 276 -413 280
rect -409 276 -407 280
rect -405 292 -404 296
rect -405 276 -400 292
rect -375 292 -374 296
rect -492 272 -452 273
rect -492 268 -456 272
rect -511 238 -510 242
rect -536 220 -531 236
rect -532 216 -531 220
rect -529 232 -528 236
rect -529 216 -524 232
rect -515 222 -510 238
rect -508 226 -500 242
rect -508 222 -506 226
rect -502 222 -500 226
rect -498 238 -497 242
rect -498 222 -493 238
rect -464 212 -459 248
rect -460 208 -459 212
rect -457 208 -449 248
rect -447 244 -446 248
rect -447 208 -442 244
rect -379 256 -374 292
rect -372 256 -364 296
rect -362 260 -357 296
rect -223 289 -218 325
rect -216 289 -208 329
rect -206 293 -201 329
rect -168 319 -167 323
rect -172 303 -167 319
rect -165 307 -157 323
rect -165 303 -163 307
rect -159 303 -157 307
rect -155 319 -154 323
rect -155 303 -150 319
rect -137 313 -136 317
rect -206 289 -205 293
rect -362 256 -361 260
rect -347 270 -346 274
rect -351 254 -346 270
rect -344 258 -339 274
rect -141 297 -136 313
rect -134 301 -129 317
rect -134 297 -133 301
rect -344 254 -343 258
rect -116 225 -111 241
rect -112 221 -111 225
rect -109 237 -108 241
rect -109 221 -104 237
rect -98 227 -93 263
rect -94 223 -93 227
rect -91 223 -83 263
rect -81 259 -80 263
rect -81 223 -76 259
rect 6 249 7 253
rect -60 239 -59 243
rect -64 223 -59 239
rect -57 227 -49 243
rect -57 223 -55 227
rect -51 223 -49 227
rect -47 239 -46 243
rect -47 223 -42 239
rect -29 233 -28 237
rect -397 184 -392 200
rect -393 180 -392 184
rect -390 186 -383 200
rect -390 182 -388 186
rect -384 182 -383 186
rect -390 180 -383 182
rect -381 196 -380 200
rect -381 180 -376 196
rect -356 196 -355 200
rect -360 180 -355 196
rect -353 184 -348 200
rect -33 217 -28 233
rect -26 221 -21 237
rect -26 217 -25 221
rect 2 213 7 249
rect 9 213 17 253
rect 19 217 24 253
rect 19 213 20 217
rect 34 227 35 231
rect -353 180 -352 184
rect -290 185 -289 189
rect -653 173 -652 177
rect -657 157 -652 173
rect -650 161 -645 177
rect -650 157 -649 161
rect -629 173 -628 177
rect -728 120 -723 136
rect -724 116 -723 120
rect -721 122 -714 136
rect -721 118 -719 122
rect -715 118 -714 122
rect -721 116 -714 118
rect -712 132 -711 136
rect -712 116 -707 132
rect -687 132 -686 136
rect -691 116 -686 132
rect -684 120 -679 136
rect -633 137 -628 173
rect -626 137 -618 177
rect -616 141 -611 177
rect -616 137 -615 141
rect -601 151 -600 155
rect -684 116 -683 120
rect -605 135 -600 151
rect -598 139 -593 155
rect -598 135 -597 139
rect -580 151 -579 155
rect -584 135 -579 151
rect -577 139 -569 155
rect -577 135 -575 139
rect -571 135 -569 139
rect -567 151 -566 155
rect -567 135 -562 151
rect -315 167 -310 183
rect -311 163 -310 167
rect -308 179 -307 183
rect -308 163 -303 179
rect -294 169 -289 185
rect -287 173 -279 189
rect -287 169 -285 173
rect -281 169 -279 173
rect -277 185 -276 189
rect -277 169 -272 185
rect -257 158 -252 194
rect -253 154 -252 158
rect -250 154 -242 194
rect -240 190 -239 194
rect -240 154 -235 190
rect 30 211 35 227
rect 37 215 42 231
rect 37 211 38 215
rect 65 227 66 231
rect 61 211 66 227
rect 68 215 76 231
rect 68 211 70 215
rect 74 211 76 215
rect 78 227 79 231
rect 78 211 83 227
rect -534 132 -529 148
rect -530 128 -529 132
rect -527 134 -520 148
rect -527 130 -525 134
rect -521 130 -520 134
rect -527 128 -520 130
rect -518 144 -517 148
rect -518 128 -513 144
rect -493 144 -492 148
rect -497 128 -492 144
rect -490 132 -485 148
rect -490 128 -489 132
rect -202 142 -197 158
rect -198 138 -197 142
rect -195 154 -194 158
rect -195 138 -190 154
rect -170 154 -169 158
rect -174 138 -169 154
rect -167 144 -160 158
rect -167 140 -166 144
rect -162 140 -160 144
rect -167 138 -160 140
rect -158 142 -153 158
rect -13 157 23 161
rect -17 156 23 157
rect -17 146 23 154
rect -158 138 -157 142
rect -17 143 23 144
rect -17 139 19 143
rect -65 114 -64 118
rect -69 98 -64 114
rect -62 102 -54 118
rect -62 98 -60 102
rect -56 98 -54 102
rect -52 114 -51 118
rect -52 98 -47 114
rect -31 114 -30 118
rect -35 98 -30 114
rect -28 102 -20 118
rect -28 98 -26 102
rect -22 98 -20 102
rect -18 114 -17 118
rect -18 98 -13 114
rect -678 45 -677 49
rect -682 29 -677 45
rect -675 47 -668 49
rect -675 43 -673 47
rect -669 43 -668 47
rect -675 29 -668 43
rect -666 33 -661 49
rect -666 29 -665 33
rect -645 33 -640 49
rect -641 29 -640 33
rect -638 45 -637 49
rect -638 29 -633 45
rect -618 12 -613 48
rect -614 8 -613 12
rect -611 8 -603 48
rect -601 44 -600 48
rect -601 8 -596 44
rect -518 45 -517 49
rect -584 21 -579 37
rect -580 17 -579 21
rect -577 33 -575 37
rect -571 33 -569 37
rect -577 17 -569 33
rect -567 21 -562 37
rect -522 29 -517 45
rect -515 47 -508 49
rect -515 43 -513 47
rect -509 43 -508 47
rect -515 29 -508 43
rect -506 33 -501 49
rect -506 29 -505 33
rect -485 33 -480 49
rect -481 29 -480 33
rect -478 45 -477 49
rect -478 29 -473 45
rect -567 17 -566 21
rect -458 12 -453 48
rect -454 8 -453 12
rect -451 8 -443 48
rect -441 44 -440 48
rect -441 8 -436 44
rect -369 48 -368 52
rect -424 21 -419 37
rect -420 17 -419 21
rect -417 33 -415 37
rect -411 33 -409 37
rect -417 17 -409 33
rect -407 21 -402 37
rect -373 32 -368 48
rect -366 50 -359 52
rect -366 46 -364 50
rect -360 46 -359 50
rect -366 32 -359 46
rect -357 36 -352 52
rect -357 32 -356 36
rect -336 36 -331 52
rect -332 32 -331 36
rect -329 48 -328 52
rect -329 32 -324 48
rect -407 17 -406 21
rect -309 15 -304 51
rect -305 11 -304 15
rect -302 11 -294 51
rect -292 47 -291 51
rect -292 11 -287 47
rect -217 48 -216 52
rect -275 24 -270 40
rect -271 20 -270 24
rect -268 36 -266 40
rect -262 36 -260 40
rect -268 20 -260 36
rect -258 24 -253 40
rect -221 32 -216 48
rect -214 50 -207 52
rect -214 46 -212 50
rect -208 46 -207 50
rect -214 32 -207 46
rect -205 36 -200 52
rect -205 32 -204 36
rect -184 36 -179 52
rect -180 32 -179 36
rect -177 48 -176 52
rect -177 32 -172 48
rect -258 20 -257 24
rect -157 15 -152 51
rect -153 11 -152 15
rect -150 11 -142 51
rect -140 47 -139 51
rect -140 11 -135 47
rect -123 24 -118 40
rect -119 20 -118 24
rect -116 36 -114 40
rect -110 36 -108 40
rect -116 20 -108 36
rect -106 24 -101 40
rect -106 20 -105 24
<< ndcontact >>
rect -159 385 -155 389
rect -153 377 -149 381
rect -149 367 -145 371
rect -155 358 -151 362
rect -149 349 -145 353
rect -326 319 -322 323
rect -265 335 -261 339
rect -247 319 -243 323
rect -318 313 -314 317
rect -308 309 -304 313
rect -299 315 -295 319
rect -290 309 -286 313
rect -510 304 -506 308
rect -516 296 -512 300
rect -520 286 -516 290
rect -514 277 -510 281
rect -520 268 -516 272
rect -422 238 -418 242
rect -404 254 -400 258
rect -223 261 -219 265
rect -214 267 -210 271
rect -172 265 -168 269
rect -154 281 -150 285
rect -141 275 -137 279
rect -133 281 -129 285
rect -205 261 -201 265
rect -379 228 -375 232
rect -370 234 -366 238
rect -351 232 -347 236
rect -343 238 -339 242
rect -361 228 -357 232
rect -536 200 -532 204
rect -528 194 -524 198
rect -515 200 -511 204
rect -116 205 -112 209
rect -497 184 -493 188
rect -464 180 -460 184
rect -455 186 -451 190
rect -446 180 -442 184
rect -108 199 -104 203
rect -98 195 -94 199
rect -89 201 -85 205
rect -80 195 -76 199
rect -657 135 -653 139
rect -649 141 -645 145
rect -397 163 -393 167
rect -388 163 -384 167
rect -380 157 -376 161
rect -360 158 -356 162
rect -352 158 -348 162
rect -64 185 -60 189
rect -46 201 -42 205
rect -33 195 -29 199
rect -25 201 -21 205
rect 2 185 6 189
rect 11 191 15 195
rect 30 189 34 193
rect 38 195 42 199
rect 20 185 24 189
rect 61 173 65 177
rect 79 189 83 193
rect -633 109 -629 113
rect -624 115 -620 119
rect -605 113 -601 117
rect -597 119 -593 123
rect -315 147 -311 151
rect -307 141 -303 145
rect -294 147 -290 151
rect 47 157 51 161
rect 41 148 45 152
rect 47 139 51 143
rect -276 131 -272 135
rect -615 109 -611 113
rect -728 99 -724 103
rect -719 99 -715 103
rect -711 93 -707 97
rect -691 94 -687 98
rect -683 94 -679 98
rect -584 97 -580 101
rect -566 113 -562 117
rect -257 126 -253 130
rect -248 132 -244 136
rect -239 126 -235 130
rect -202 116 -198 120
rect -194 116 -190 120
rect -534 111 -530 115
rect -525 111 -521 115
rect -517 105 -513 109
rect -497 106 -493 110
rect -174 115 -170 119
rect -166 121 -162 125
rect -157 121 -153 125
rect -489 106 -485 110
rect -682 62 -678 66
rect -673 62 -669 66
rect -665 68 -661 72
rect -618 72 -614 76
rect -645 67 -641 71
rect -637 67 -633 71
rect -609 66 -605 70
rect -600 72 -596 76
rect -584 71 -580 75
rect -522 62 -518 66
rect -513 62 -509 66
rect -505 68 -501 72
rect -458 72 -454 76
rect -485 67 -481 71
rect -566 55 -562 59
rect -477 67 -473 71
rect -449 66 -445 70
rect -440 72 -436 76
rect -424 71 -420 75
rect -373 65 -369 69
rect -364 65 -360 69
rect -356 71 -352 75
rect -309 75 -305 79
rect -336 70 -332 74
rect -406 55 -402 59
rect -328 70 -324 74
rect -300 69 -296 73
rect -291 75 -287 79
rect -275 74 -271 78
rect -221 65 -217 69
rect -212 65 -208 69
rect -204 71 -200 75
rect -157 75 -153 79
rect -184 70 -180 74
rect -257 58 -253 62
rect -176 70 -172 74
rect -148 69 -144 73
rect -139 75 -135 79
rect -123 74 -119 78
rect -105 58 -101 62
rect -69 60 -65 64
rect -51 76 -47 80
rect -35 60 -31 64
rect -17 76 -13 80
<< pdcontact >>
rect -175 385 -171 389
rect -191 377 -187 381
rect -326 335 -322 339
rect -318 351 -314 355
rect -308 337 -304 341
rect -290 373 -286 377
rect -265 373 -261 377
rect -256 357 -252 361
rect -247 373 -243 377
rect -177 367 -173 371
rect -213 349 -209 353
rect -223 325 -219 329
rect -494 304 -490 308
rect -478 296 -474 300
rect -422 292 -418 296
rect -492 286 -488 290
rect -413 276 -409 280
rect -404 292 -400 296
rect -379 292 -375 296
rect -456 268 -452 272
rect -515 238 -511 242
rect -536 216 -532 220
rect -528 232 -524 236
rect -506 222 -502 226
rect -497 238 -493 242
rect -464 208 -460 212
rect -446 244 -442 248
rect -172 319 -168 323
rect -163 303 -159 307
rect -154 319 -150 323
rect -141 313 -137 317
rect -205 289 -201 293
rect -361 256 -357 260
rect -351 270 -347 274
rect -133 297 -129 301
rect -343 254 -339 258
rect -116 221 -112 225
rect -108 237 -104 241
rect -98 223 -94 227
rect -80 259 -76 263
rect 2 249 6 253
rect -64 239 -60 243
rect -55 223 -51 227
rect -46 239 -42 243
rect -33 233 -29 237
rect -397 180 -393 184
rect -388 182 -384 186
rect -380 196 -376 200
rect -360 196 -356 200
rect -25 217 -21 221
rect 20 213 24 217
rect 30 227 34 231
rect -352 180 -348 184
rect -294 185 -290 189
rect -657 173 -653 177
rect -649 157 -645 161
rect -633 173 -629 177
rect -728 116 -724 120
rect -719 118 -715 122
rect -711 132 -707 136
rect -691 132 -687 136
rect -615 137 -611 141
rect -605 151 -601 155
rect -683 116 -679 120
rect -597 135 -593 139
rect -584 151 -580 155
rect -575 135 -571 139
rect -566 151 -562 155
rect -315 163 -311 167
rect -307 179 -303 183
rect -285 169 -281 173
rect -276 185 -272 189
rect -257 154 -253 158
rect -239 190 -235 194
rect 38 211 42 215
rect 61 227 65 231
rect 70 211 74 215
rect 79 227 83 231
rect -534 128 -530 132
rect -525 130 -521 134
rect -517 144 -513 148
rect -497 144 -493 148
rect -489 128 -485 132
rect -202 138 -198 142
rect -194 154 -190 158
rect -174 154 -170 158
rect -166 140 -162 144
rect -17 157 -13 161
rect -157 138 -153 142
rect 19 139 23 143
rect -69 114 -65 118
rect -60 98 -56 102
rect -51 114 -47 118
rect -35 114 -31 118
rect -26 98 -22 102
rect -17 114 -13 118
rect -682 45 -678 49
rect -673 43 -669 47
rect -665 29 -661 33
rect -645 29 -641 33
rect -637 45 -633 49
rect -618 8 -614 12
rect -600 44 -596 48
rect -522 45 -518 49
rect -584 17 -580 21
rect -575 33 -571 37
rect -513 43 -509 47
rect -505 29 -501 33
rect -485 29 -481 33
rect -477 45 -473 49
rect -566 17 -562 21
rect -458 8 -454 12
rect -440 44 -436 48
rect -373 48 -369 52
rect -424 17 -420 21
rect -415 33 -411 37
rect -364 46 -360 50
rect -356 32 -352 36
rect -336 32 -332 36
rect -328 48 -324 52
rect -406 17 -402 21
rect -309 11 -305 15
rect -291 47 -287 51
rect -221 48 -217 52
rect -275 20 -271 24
rect -266 36 -262 40
rect -212 46 -208 50
rect -204 32 -200 36
rect -184 32 -180 36
rect -176 48 -172 52
rect -257 20 -253 24
rect -157 11 -153 15
rect -139 47 -135 51
rect -123 20 -119 24
rect -114 36 -110 40
rect -105 20 -101 24
<< polysilicon >>
rect -194 382 -191 384
rect -171 382 -159 384
rect -149 382 -146 384
rect -303 377 -301 380
rect -293 377 -291 380
rect -260 377 -258 381
rect -250 377 -248 381
rect -321 355 -319 358
rect -216 364 -213 366
rect -173 364 -155 366
rect -145 364 -142 366
rect -260 339 -258 357
rect -250 339 -248 357
rect -216 354 -213 356
rect -173 354 -155 356
rect -145 354 -142 356
rect -321 323 -319 335
rect -303 319 -301 337
rect -293 319 -291 337
rect -218 329 -216 332
rect -208 329 -206 332
rect -321 310 -319 313
rect -260 315 -258 319
rect -250 315 -248 319
rect -303 306 -301 309
rect -293 306 -291 309
rect -519 301 -516 303
rect -506 301 -494 303
rect -474 301 -471 303
rect -417 296 -415 300
rect -407 296 -405 300
rect -374 296 -372 299
rect -364 296 -362 299
rect -523 283 -520 285
rect -510 283 -492 285
rect -452 283 -449 285
rect -523 273 -520 275
rect -510 273 -492 275
rect -452 273 -449 275
rect -417 258 -415 276
rect -407 258 -405 276
rect -459 248 -457 251
rect -449 248 -447 251
rect -510 242 -508 246
rect -500 242 -498 246
rect -531 236 -529 240
rect -531 204 -529 216
rect -510 204 -508 222
rect -500 204 -498 222
rect -167 323 -165 327
rect -157 323 -155 327
rect -136 317 -134 321
rect -346 274 -344 277
rect -374 238 -372 256
rect -364 238 -362 256
rect -218 271 -216 289
rect -208 271 -206 289
rect -167 285 -165 303
rect -157 285 -155 303
rect -136 285 -134 297
rect -136 271 -134 275
rect -167 261 -165 265
rect -157 261 -155 265
rect -93 263 -91 266
rect -83 263 -81 266
rect -218 258 -216 261
rect -208 258 -206 261
rect -346 242 -344 254
rect -417 234 -415 238
rect -407 234 -405 238
rect -111 241 -109 244
rect -346 229 -344 232
rect -374 225 -372 228
rect -364 225 -362 228
rect 7 253 9 256
rect 17 253 19 256
rect -59 243 -57 247
rect -49 243 -47 247
rect -28 237 -26 241
rect -531 190 -529 194
rect -459 190 -457 208
rect -449 190 -447 208
rect -392 200 -390 212
rect -111 209 -109 221
rect -383 200 -381 203
rect -355 200 -353 204
rect -652 177 -650 181
rect -510 180 -508 184
rect -500 180 -498 184
rect -93 205 -91 223
rect -83 205 -81 223
rect -59 205 -57 223
rect -49 205 -47 223
rect -28 205 -26 217
rect 35 231 37 234
rect 66 231 68 235
rect 76 231 78 235
rect -252 194 -250 197
rect -242 194 -240 197
rect -111 196 -109 199
rect -289 189 -287 193
rect -279 189 -277 193
rect -310 183 -308 187
rect -628 177 -626 180
rect -618 177 -616 180
rect -459 177 -457 180
rect -449 177 -447 180
rect -723 136 -721 148
rect -652 145 -650 157
rect -714 136 -712 139
rect -686 136 -684 140
rect -392 174 -390 180
rect -392 167 -390 171
rect -383 167 -381 180
rect -355 168 -353 180
rect -600 155 -598 158
rect -579 155 -577 159
rect -569 155 -567 159
rect -652 131 -650 135
rect -628 119 -626 137
rect -618 119 -616 137
rect -529 148 -527 160
rect -392 155 -390 157
rect -520 148 -518 151
rect -492 148 -490 152
rect -392 151 -391 155
rect -383 154 -381 157
rect -355 154 -353 158
rect -310 151 -308 163
rect -289 151 -287 169
rect -279 151 -277 169
rect -93 192 -91 195
rect -83 192 -81 195
rect 7 195 9 213
rect 17 195 19 213
rect 35 199 37 211
rect -28 191 -26 195
rect 66 193 68 211
rect 76 193 78 211
rect 35 186 37 189
rect -59 181 -57 185
rect -49 181 -47 185
rect 7 182 9 185
rect 17 182 19 185
rect -197 158 -195 162
rect -169 158 -167 161
rect -160 158 -158 170
rect 66 169 68 173
rect 76 169 78 173
rect -392 150 -390 151
rect -600 123 -598 135
rect -723 110 -721 116
rect -723 103 -721 107
rect -714 103 -712 116
rect -686 104 -684 116
rect -579 117 -577 135
rect -569 117 -567 135
rect -310 137 -308 141
rect -252 136 -250 154
rect -242 136 -240 154
rect -20 154 -17 156
rect 23 154 41 156
rect 51 154 54 156
rect -20 144 -17 146
rect 23 144 41 146
rect 51 144 54 146
rect -529 122 -527 128
rect -600 110 -598 113
rect -628 106 -626 109
rect -618 106 -616 109
rect -529 115 -527 119
rect -520 115 -518 128
rect -492 116 -490 128
rect -289 127 -287 131
rect -279 127 -277 131
rect -197 126 -195 138
rect -252 123 -250 126
rect -242 123 -240 126
rect -169 125 -167 138
rect -160 132 -158 138
rect -160 125 -158 129
rect -197 112 -195 116
rect -64 118 -62 122
rect -54 118 -52 122
rect -30 118 -28 122
rect -20 118 -18 122
rect -169 112 -167 115
rect -160 113 -158 115
rect -159 109 -158 113
rect -160 108 -158 109
rect -529 103 -527 105
rect -529 99 -528 103
rect -520 102 -518 105
rect -492 102 -490 106
rect -529 98 -527 99
rect -723 91 -721 93
rect -723 87 -722 91
rect -714 90 -712 93
rect -686 90 -684 94
rect -579 93 -577 97
rect -569 93 -567 97
rect -723 86 -721 87
rect -368 81 -366 82
rect -677 78 -675 79
rect -677 74 -676 78
rect -613 76 -611 79
rect -603 76 -601 79
rect -677 72 -675 74
rect -668 72 -666 75
rect -640 71 -638 75
rect -677 58 -675 62
rect -677 49 -675 55
rect -668 49 -666 62
rect -579 75 -577 79
rect -569 75 -567 79
rect -517 78 -515 79
rect -640 49 -638 61
rect -613 48 -611 66
rect -603 48 -601 66
rect -517 74 -516 78
rect -453 76 -451 79
rect -443 76 -441 79
rect -517 72 -515 74
rect -508 72 -506 75
rect -480 71 -478 75
rect -517 58 -515 62
rect -677 17 -675 29
rect -668 26 -666 29
rect -640 25 -638 29
rect -579 37 -577 55
rect -569 37 -567 55
rect -517 49 -515 55
rect -508 49 -506 62
rect -419 75 -417 79
rect -409 75 -407 79
rect -368 77 -367 81
rect -304 79 -302 82
rect -294 79 -292 82
rect -368 75 -366 77
rect -359 75 -357 78
rect -480 49 -478 61
rect -453 48 -451 66
rect -443 48 -441 66
rect -331 74 -329 78
rect -368 61 -366 65
rect -517 17 -515 29
rect -508 26 -506 29
rect -480 25 -478 29
rect -579 13 -577 17
rect -569 13 -567 17
rect -419 37 -417 55
rect -409 37 -407 55
rect -368 52 -366 58
rect -359 52 -357 65
rect -270 78 -268 82
rect -260 78 -258 82
rect -216 81 -214 82
rect -331 52 -329 64
rect -304 51 -302 69
rect -294 51 -292 69
rect -216 77 -215 81
rect -152 79 -150 82
rect -142 79 -140 82
rect -216 75 -214 77
rect -207 75 -205 78
rect -179 74 -177 78
rect -216 61 -214 65
rect -368 20 -366 32
rect -359 29 -357 32
rect -331 28 -329 32
rect -419 13 -417 17
rect -409 13 -407 17
rect -270 40 -268 58
rect -260 40 -258 58
rect -216 52 -214 58
rect -207 52 -205 65
rect -118 78 -116 82
rect -108 78 -106 82
rect -64 80 -62 98
rect -54 80 -52 98
rect -30 80 -28 98
rect -20 80 -18 98
rect -179 52 -177 64
rect -152 51 -150 69
rect -142 51 -140 69
rect -216 20 -214 32
rect -207 29 -205 32
rect -179 28 -177 32
rect -270 16 -268 20
rect -260 16 -258 20
rect -118 40 -116 58
rect -108 40 -106 58
rect -64 56 -62 60
rect -54 56 -52 60
rect -30 56 -28 60
rect -20 56 -18 60
rect -118 16 -116 20
rect -108 16 -106 20
rect -304 8 -302 11
rect -294 8 -292 11
rect -152 8 -150 11
rect -142 8 -140 11
rect -613 5 -611 8
rect -603 5 -601 8
rect -453 5 -451 8
rect -443 5 -441 8
<< polycontact >>
rect -164 378 -160 382
rect -258 340 -254 344
rect -166 360 -162 364
rect -248 346 -244 350
rect -160 350 -156 354
rect -319 324 -315 328
rect -301 326 -297 330
rect -291 320 -287 324
rect -505 297 -501 301
rect -503 279 -499 283
rect -509 269 -505 273
rect -421 265 -417 269
rect -411 259 -407 263
rect -529 205 -525 209
rect -508 205 -504 209
rect -498 211 -494 215
rect -171 292 -167 296
rect -378 239 -374 243
rect -368 245 -364 249
rect -222 272 -218 276
rect -212 278 -208 282
rect -161 286 -157 290
rect -140 286 -136 290
rect -350 243 -346 247
rect -457 197 -453 201
rect -390 207 -386 211
rect -109 210 -105 214
rect -447 191 -443 195
rect -91 212 -87 216
rect -63 213 -59 217
rect -81 206 -77 210
rect -53 206 -49 210
rect -32 206 -28 210
rect -721 143 -717 147
rect -656 146 -652 150
rect -381 169 -377 173
rect -359 169 -355 173
rect -632 120 -628 124
rect -622 126 -618 130
rect -527 155 -523 159
rect -391 151 -387 155
rect -308 152 -304 156
rect -287 152 -283 156
rect -277 158 -273 162
rect 3 196 7 200
rect 13 202 17 206
rect 31 200 35 204
rect 62 200 66 204
rect 72 194 76 198
rect -164 165 -160 169
rect -604 124 -600 128
rect -583 124 -579 128
rect -712 105 -708 109
rect -690 105 -686 109
rect -573 118 -569 122
rect -250 143 -246 147
rect -240 137 -236 141
rect 36 156 40 160
rect 30 146 34 150
rect -518 117 -514 121
rect -496 117 -492 121
rect -195 127 -191 131
rect -173 127 -169 131
rect -163 109 -159 113
rect -528 99 -524 103
rect -722 87 -718 91
rect -68 87 -64 91
rect -676 74 -672 78
rect -617 61 -613 65
rect -666 56 -662 60
rect -644 56 -640 60
rect -607 55 -603 59
rect -516 74 -512 78
rect -675 18 -671 22
rect -583 44 -579 48
rect -573 50 -569 54
rect -367 77 -363 81
rect -457 61 -453 65
rect -506 56 -502 60
rect -484 56 -480 60
rect -447 55 -443 59
rect -515 18 -511 22
rect -423 44 -419 48
rect -413 50 -409 54
rect -308 64 -304 68
rect -357 59 -353 63
rect -335 59 -331 63
rect -298 58 -294 62
rect -215 77 -211 81
rect -366 21 -362 25
rect -274 47 -270 51
rect -264 53 -260 57
rect -58 81 -54 85
rect -34 87 -30 91
rect -24 81 -20 85
rect -156 64 -152 68
rect -205 59 -201 63
rect -183 59 -179 63
rect -146 58 -142 62
rect -214 21 -210 25
rect -122 47 -118 51
rect -112 53 -108 57
<< metal1 >>
rect -201 393 -161 396
rect -317 384 -242 387
rect -201 387 -198 393
rect -164 389 -161 393
rect -229 384 -198 387
rect -171 386 -159 389
rect -317 366 -314 384
rect -289 377 -286 384
rect -265 377 -261 384
rect -246 377 -243 384
rect -341 363 -314 366
rect -504 312 -464 315
rect -504 308 -501 312
rect -506 305 -494 308
rect -467 306 -464 312
rect -467 303 -436 306
rect -341 306 -338 363
rect -317 355 -314 363
rect -256 356 -253 357
rect -265 353 -253 356
rect -265 344 -262 353
rect -229 350 -226 384
rect -244 347 -226 350
rect -218 377 -191 380
rect -223 352 -220 375
rect -164 371 -161 378
rect -149 377 -138 380
rect -141 371 -138 377
rect -173 368 -156 371
rect -159 362 -156 368
rect -145 368 -138 371
rect -223 349 -213 352
rect -283 341 -262 344
rect -326 328 -323 335
rect -308 328 -305 337
rect -283 330 -280 341
rect -265 339 -262 341
rect -254 340 -235 343
rect -238 337 -235 340
rect -223 339 -220 349
rect -166 343 -163 360
rect -159 359 -155 362
rect -141 353 -138 368
rect -160 348 -156 350
rect -145 349 -141 352
rect -160 346 -159 348
rect -223 336 -175 339
rect -132 341 -129 451
rect -132 338 -106 341
rect -328 323 -323 328
rect -315 325 -305 328
rect -297 327 -280 330
rect -223 329 -220 336
rect -178 333 -175 336
rect -178 330 -114 333
rect -308 323 -305 325
rect -308 320 -296 323
rect -287 321 -283 324
rect -299 319 -296 320
rect -172 323 -169 330
rect -154 323 -150 330
rect -246 314 -243 319
rect -141 317 -138 330
rect -423 303 -338 306
rect -317 305 -314 313
rect -308 305 -305 309
rect -289 305 -286 309
rect -282 311 -234 314
rect -282 305 -279 311
rect -527 296 -516 299
rect -527 290 -524 296
rect -504 290 -501 297
rect -474 296 -447 299
rect -527 287 -520 290
rect -527 272 -524 287
rect -509 287 -492 290
rect -509 281 -506 287
rect -510 278 -506 281
rect -524 268 -520 271
rect -508 264 -505 269
rect -556 260 -505 264
rect -502 262 -499 279
rect -445 271 -442 294
rect -452 268 -442 271
rect -445 258 -442 268
rect -439 269 -436 303
rect -422 296 -419 303
rect -404 296 -400 303
rect -379 296 -376 303
rect -412 275 -409 276
rect -412 272 -400 275
rect -439 266 -421 269
rect -403 263 -400 272
rect -351 274 -348 303
rect -326 302 -279 305
rect -490 255 -442 258
rect -425 259 -411 262
rect -403 260 -382 263
rect -403 258 -400 260
rect -490 252 -487 255
rect -566 249 -487 252
rect -673 186 -602 187
rect -673 184 -590 186
rect -673 183 -663 184
rect -673 156 -669 183
rect -657 177 -654 184
rect -633 177 -630 184
rect -605 183 -590 184
rect -605 165 -602 183
rect -593 176 -590 183
rect -566 176 -563 249
rect -527 236 -524 249
rect -515 242 -511 249
rect -496 242 -493 249
rect -445 248 -442 255
rect -385 249 -382 260
rect -385 246 -368 249
rect -360 247 -357 256
rect -342 247 -339 254
rect -360 244 -350 247
rect -382 240 -378 243
rect -360 242 -357 244
rect -342 244 -336 247
rect -342 242 -339 244
rect -369 239 -357 242
rect -369 238 -366 239
rect -422 233 -419 238
rect -431 230 -383 233
rect -506 221 -503 222
rect -515 218 -503 221
rect -536 209 -533 216
rect -515 209 -512 218
rect -494 212 -467 215
rect -539 206 -533 209
rect -536 204 -533 206
rect -525 206 -512 209
rect -515 204 -512 206
rect -504 205 -490 208
rect -470 199 -467 212
rect -464 199 -461 208
rect -470 196 -461 199
rect -453 198 -440 201
rect -527 180 -524 194
rect -464 194 -461 196
rect -464 191 -452 194
rect -443 192 -435 195
rect -455 190 -452 191
rect -530 177 -528 180
rect -593 173 -563 176
rect -496 179 -493 184
rect -523 176 -487 179
rect -464 176 -461 180
rect -445 176 -442 180
rect -431 176 -428 230
rect -386 224 -383 230
rect -379 224 -376 228
rect -360 224 -357 228
rect -351 224 -348 232
rect -326 224 -323 302
rect -237 257 -234 311
rect -162 302 -159 303
rect -162 299 -150 302
rect -198 293 -171 296
rect -225 279 -212 282
rect -204 280 -201 289
rect -198 280 -195 293
rect -153 290 -150 299
rect -132 290 -129 297
rect -185 286 -161 289
rect -153 287 -140 290
rect -185 284 -181 286
rect -153 285 -150 287
rect -132 287 -126 290
rect -132 285 -129 287
rect -204 277 -195 280
rect -231 275 -222 276
rect -226 273 -222 275
rect -204 275 -201 277
rect -213 272 -201 275
rect -213 271 -210 272
rect -223 257 -220 261
rect -204 257 -201 261
rect -172 260 -169 265
rect -141 261 -138 275
rect -117 273 -114 330
rect -109 282 -106 338
rect -109 279 -59 282
rect -117 270 -66 273
rect -178 257 -142 260
rect -237 254 -174 257
rect -107 251 -104 270
rect -79 263 -76 270
rect -118 248 -104 251
rect -69 253 -66 270
rect -62 271 -59 279
rect -62 268 41 271
rect -33 260 33 263
rect -33 253 -30 260
rect -69 250 -30 253
rect -107 241 -104 248
rect -64 243 -61 250
rect -46 243 -42 250
rect -33 237 -30 250
rect 2 253 5 260
rect 30 241 33 260
rect 38 248 41 268
rect 38 245 101 248
rect 30 238 89 241
rect 30 231 33 238
rect 61 231 64 238
rect 79 231 83 238
rect -386 221 -323 224
rect -116 214 -113 221
rect -98 214 -95 223
rect -54 222 -51 223
rect -54 219 -42 222
rect -386 208 -375 210
rect -123 211 -113 214
rect -116 209 -113 211
rect -105 211 -95 214
rect -87 213 -63 216
rect -98 209 -95 211
rect -45 210 -42 219
rect -24 210 -21 217
rect -386 207 -371 208
rect -374 200 -371 207
rect -360 205 -342 209
rect -98 206 -86 209
rect -77 207 -53 210
rect -45 207 -32 210
rect -89 205 -86 206
rect -45 205 -42 207
rect -24 205 -17 210
rect -360 200 -356 205
rect -376 197 -363 200
rect -491 173 -428 176
rect -396 173 -393 180
rect -388 179 -385 182
rect -561 165 -493 168
rect -605 162 -556 165
rect -746 152 -669 156
rect -746 79 -742 152
rect -717 143 -702 146
rect -705 136 -702 143
rect -691 136 -687 152
rect -648 150 -645 157
rect -605 155 -602 162
rect -584 155 -581 162
rect -566 155 -562 162
rect -497 160 -493 165
rect -511 158 -508 160
rect -523 155 -508 158
rect -511 152 -508 155
rect -497 157 -478 160
rect -660 147 -656 150
rect -648 147 -637 150
rect -511 148 -510 152
rect -648 145 -645 147
rect -707 133 -694 136
rect -727 109 -724 116
rect -719 115 -716 118
rect -736 107 -724 109
rect -731 106 -724 107
rect -727 103 -724 106
rect -719 103 -716 110
rect -697 109 -694 133
rect -708 105 -705 108
rect -697 106 -690 109
rect -707 92 -701 96
rect -707 90 -706 92
rect -718 87 -706 90
rect -746 75 -704 79
rect -697 78 -694 106
rect -682 100 -679 116
rect -682 98 -678 100
rect -679 95 -678 98
rect -691 89 -688 94
rect -657 89 -654 135
rect -640 130 -637 147
rect -513 147 -510 148
rect -497 148 -493 157
rect -505 147 -500 148
rect -513 145 -500 147
rect -640 127 -622 130
rect -614 128 -611 137
rect -596 128 -593 135
rect -574 134 -571 135
rect -574 131 -562 134
rect -614 125 -604 128
rect -635 121 -632 124
rect -614 123 -611 125
rect -596 125 -583 128
rect -596 123 -593 125
rect -623 120 -611 123
rect -623 119 -620 120
rect -565 122 -562 131
rect -585 118 -573 121
rect -565 121 -542 122
rect -533 121 -530 128
rect -525 127 -522 130
rect -565 119 -530 121
rect -565 117 -562 119
rect -633 105 -630 109
rect -614 105 -611 109
rect -605 106 -602 113
rect -558 109 -555 119
rect -545 118 -542 119
rect -537 118 -530 119
rect -533 115 -530 118
rect -525 115 -522 122
rect -503 121 -500 145
rect -514 117 -511 120
rect -503 118 -496 121
rect -488 112 -485 128
rect -488 110 -484 112
rect -644 102 -606 105
rect -644 89 -641 102
rect -513 104 -507 108
rect -513 102 -512 104
rect -524 99 -512 102
rect -485 107 -484 110
rect -497 101 -494 106
rect -475 101 -472 173
rect -408 171 -393 173
rect -408 170 -405 171
rect -400 170 -393 171
rect -396 167 -393 170
rect -388 167 -385 174
rect -366 173 -363 197
rect -346 200 -342 205
rect -269 201 -217 204
rect -346 199 -302 200
rect -269 199 -266 201
rect -346 196 -266 199
rect -306 183 -303 196
rect -294 189 -290 196
rect -275 189 -272 196
rect -238 194 -235 201
rect -377 169 -374 172
rect -366 170 -359 173
rect -351 164 -348 180
rect -220 170 -217 201
rect -21 201 -17 205
rect 0 203 13 206
rect 21 204 24 213
rect 39 204 42 211
rect 71 210 74 211
rect 71 207 83 210
rect -107 191 -104 199
rect -98 191 -95 195
rect -79 191 -76 195
rect -129 188 -68 191
rect -285 168 -282 169
rect -351 162 -347 164
rect -376 156 -370 160
rect -376 154 -375 156
rect -387 151 -375 154
rect -348 159 -347 162
rect -294 165 -282 168
rect -220 167 -190 170
rect -360 153 -357 158
rect -315 156 -312 163
rect -294 156 -291 165
rect -273 159 -266 162
rect -194 158 -190 167
rect -179 168 -176 170
rect -179 165 -164 168
rect -179 158 -176 165
rect -326 153 -312 156
rect -360 150 -355 153
rect -360 146 -357 150
rect -445 143 -357 146
rect -445 111 -442 143
rect -326 131 -323 153
rect -315 151 -312 153
rect -304 153 -291 156
rect -294 151 -291 153
rect -283 152 -266 155
rect -269 145 -266 152
rect -187 155 -174 158
rect -257 145 -254 154
rect -269 142 -254 145
rect -246 144 -221 147
rect -365 128 -323 131
rect -365 114 -362 128
rect -306 126 -303 141
rect -257 140 -254 142
rect -257 137 -245 140
rect -236 137 -234 141
rect -248 136 -245 137
rect -275 126 -272 131
rect -306 123 -266 126
rect -269 122 -266 123
rect -257 122 -254 126
rect -238 122 -235 126
rect -269 119 -228 122
rect -365 111 -351 114
rect -445 108 -379 111
rect -497 98 -472 101
rect -584 93 -581 97
rect -691 86 -641 89
rect -475 92 -472 98
rect -382 96 -379 108
rect -580 89 -472 92
rect -645 83 -641 86
rect -475 83 -472 89
rect -405 93 -333 96
rect -405 83 -402 93
rect -645 80 -581 83
rect -708 2 -704 75
rect -672 75 -660 78
rect -661 73 -660 75
rect -661 69 -655 73
rect -645 71 -642 80
rect -618 76 -615 80
rect -599 76 -596 80
rect -635 71 -632 73
rect -633 67 -632 71
rect -584 75 -581 80
rect -485 80 -402 83
rect -336 86 -333 93
rect -261 86 -258 119
rect -231 111 -228 119
rect -229 106 -228 111
rect -336 83 -253 86
rect -512 75 -500 78
rect -501 73 -500 75
rect -693 58 -690 59
rect -681 59 -678 62
rect -685 58 -678 59
rect -693 56 -678 58
rect -693 13 -690 56
rect -681 49 -678 56
rect -673 55 -670 62
rect -662 57 -659 60
rect -651 56 -644 59
rect -651 52 -648 56
rect -673 47 -670 50
rect -636 49 -633 67
rect -501 69 -495 73
rect -485 71 -482 80
rect -458 76 -455 80
rect -439 76 -436 80
rect -475 71 -472 73
rect -473 67 -472 71
rect -424 75 -421 80
rect -608 65 -605 66
rect -620 61 -617 64
rect -608 64 -596 65
rect -608 62 -593 64
rect -599 61 -588 62
rect -624 55 -607 58
rect -624 52 -621 55
rect -651 32 -648 47
rect -599 48 -596 61
rect -586 51 -573 54
rect -565 53 -562 55
rect -533 58 -530 59
rect -521 59 -518 62
rect -525 58 -518 59
rect -533 56 -518 58
rect -559 53 -556 56
rect -565 50 -556 53
rect -590 44 -583 47
rect -590 40 -587 44
rect -565 41 -562 50
rect -574 38 -562 41
rect -574 37 -571 38
rect -661 29 -648 32
rect -659 22 -656 29
rect -671 19 -656 22
rect -645 20 -641 29
rect -660 13 -657 19
rect -645 17 -621 20
rect -624 2 -621 17
rect -708 1 -621 2
rect -584 10 -581 17
rect -566 10 -562 17
rect -533 13 -530 56
rect -521 49 -518 56
rect -513 55 -510 62
rect -502 57 -499 60
rect -491 56 -484 59
rect -491 52 -488 56
rect -513 47 -510 50
rect -476 49 -473 67
rect -448 65 -445 66
rect -460 61 -457 64
rect -448 64 -436 65
rect -448 62 -433 64
rect -439 61 -428 62
rect -464 55 -447 58
rect -464 52 -461 55
rect -491 32 -488 47
rect -439 48 -436 61
rect -426 51 -413 54
rect -405 53 -402 55
rect -399 53 -396 83
rect -363 78 -351 81
rect -352 76 -351 78
rect -352 72 -346 76
rect -336 74 -333 83
rect -309 79 -306 83
rect -290 79 -287 83
rect -326 74 -323 76
rect -324 70 -323 74
rect -275 78 -272 83
rect -405 50 -396 53
rect -384 61 -381 62
rect -372 62 -369 65
rect -376 61 -369 62
rect -384 59 -369 61
rect -430 44 -423 47
rect -430 40 -427 44
rect -405 41 -402 50
rect -414 38 -402 41
rect -414 37 -411 38
rect -501 29 -488 32
rect -499 22 -496 29
rect -511 19 -496 22
rect -485 20 -481 29
rect -500 13 -497 19
rect -485 17 -461 20
rect -618 1 -615 8
rect -594 7 -556 10
rect -594 2 -590 7
rect -464 2 -461 17
rect -594 1 -461 2
rect -424 10 -421 17
rect -406 10 -402 17
rect -384 16 -381 59
rect -372 52 -369 59
rect -364 58 -361 65
rect -353 60 -350 63
rect -342 59 -335 62
rect -342 55 -339 59
rect -364 50 -361 53
rect -327 52 -324 70
rect -299 68 -296 69
rect -311 64 -308 67
rect -299 67 -287 68
rect -299 65 -284 67
rect -290 64 -279 65
rect -315 58 -298 61
rect -315 55 -312 58
rect -342 35 -339 50
rect -290 51 -287 64
rect -277 54 -264 57
rect -256 56 -253 58
rect -250 57 -247 93
rect -231 89 -228 106
rect -224 95 -221 144
rect -202 122 -199 138
rect -187 133 -184 155
rect -165 137 -162 140
rect -191 128 -190 131
rect -185 128 -184 133
rect -176 127 -173 130
rect -165 125 -162 132
rect -203 120 -199 122
rect -157 131 -154 138
rect -145 131 -142 164
rect -157 129 -142 131
rect -129 130 -126 188
rect -71 180 -68 188
rect -64 180 -61 185
rect -33 181 -30 195
rect -20 192 -17 201
rect 21 201 31 204
rect -5 198 3 199
rect 0 196 3 198
rect 21 199 24 201
rect 39 201 62 204
rect 39 199 42 201
rect 12 196 24 199
rect 12 195 15 196
rect 80 198 83 207
rect -19 187 -17 192
rect 48 194 72 197
rect 80 195 93 198
rect 48 193 52 194
rect 80 193 83 195
rect 2 181 5 185
rect 21 181 24 185
rect 30 181 33 189
rect -33 180 58 181
rect -71 178 58 180
rect -71 177 -30 178
rect -157 128 -150 129
rect -157 125 -154 128
rect -145 128 -142 129
rect -139 127 -126 130
rect -27 161 -24 163
rect -27 158 -17 161
rect -27 128 -24 158
rect 30 150 33 175
rect 55 168 58 178
rect 90 175 93 195
rect 61 168 64 173
rect 55 165 86 168
rect 36 160 39 165
rect 55 161 58 165
rect 98 161 101 245
rect 51 158 58 161
rect 37 148 41 151
rect 37 142 40 148
rect 23 139 40 142
rect 55 142 58 158
rect 51 139 58 142
rect 63 158 101 161
rect 32 131 35 139
rect 63 135 66 158
rect 15 128 35 131
rect 40 132 66 135
rect -203 117 -202 120
rect -193 111 -190 116
rect -212 108 -190 111
rect -180 114 -174 118
rect -175 112 -174 114
rect -175 109 -163 112
rect -139 102 -136 127
rect -75 125 -7 128
rect -69 118 -66 125
rect -51 118 -47 125
rect -35 118 -32 125
rect -17 118 -13 125
rect 40 124 43 132
rect 0 121 43 124
rect -139 99 -120 102
rect -224 92 -132 95
rect -231 86 -181 89
rect -123 86 -120 99
rect -59 97 -56 98
rect -25 97 -22 98
rect -59 94 -47 97
rect -25 94 -13 97
rect -184 83 -114 86
rect -211 78 -199 81
rect -200 76 -199 78
rect -200 72 -194 76
rect -184 74 -181 83
rect -157 79 -154 83
rect -138 79 -135 83
rect -174 74 -171 76
rect -172 70 -171 74
rect -123 78 -120 83
rect -232 61 -229 62
rect -220 62 -217 65
rect -224 61 -217 62
rect -232 59 -217 61
rect -256 53 -250 56
rect -281 47 -274 50
rect -281 43 -278 47
rect -256 44 -253 53
rect -265 41 -253 44
rect -265 40 -262 41
rect -352 32 -339 35
rect -350 25 -347 32
rect -362 22 -347 25
rect -336 23 -332 32
rect -351 16 -348 22
rect -336 20 -312 23
rect -315 10 -312 20
rect -458 1 -455 8
rect -434 7 -312 10
rect -434 1 -430 7
rect -315 4 -312 7
rect -275 13 -272 20
rect -257 13 -253 20
rect -232 16 -229 59
rect -220 52 -217 59
rect -212 58 -209 65
rect -201 60 -198 63
rect -190 59 -183 62
rect -190 55 -187 59
rect -212 50 -209 53
rect -175 52 -172 70
rect -147 68 -144 69
rect -159 64 -156 67
rect -147 67 -135 68
rect -147 65 -132 67
rect -138 64 -127 65
rect -163 58 -146 61
rect -163 55 -160 58
rect -190 35 -187 50
rect -138 51 -135 64
rect -125 54 -112 57
rect -104 56 -101 58
rect -98 56 -95 90
rect -74 88 -68 91
rect -104 53 -95 56
rect -82 81 -58 84
rect -50 84 -47 94
rect -36 87 -34 91
rect -16 85 -13 94
rect 0 85 3 121
rect -50 81 -24 84
rect -16 82 3 85
rect -129 47 -122 50
rect -129 43 -126 47
rect -104 44 -101 53
rect -113 41 -101 44
rect -113 40 -110 41
rect -200 32 -187 35
rect -198 25 -195 32
rect -210 22 -195 25
rect -184 23 -180 32
rect -82 29 -79 81
rect -50 80 -47 81
rect -16 80 -13 82
rect -69 56 -66 60
rect -71 55 -66 56
rect -35 55 -32 60
rect -71 52 -10 55
rect -199 16 -196 22
rect -184 20 -160 23
rect -163 13 -160 20
rect -309 4 -306 11
rect -285 10 -160 13
rect -285 4 -281 10
rect -315 1 -281 4
rect -163 4 -160 10
rect -123 13 -120 20
rect -105 13 -101 20
rect -157 4 -154 11
rect -133 10 -95 13
rect -133 4 -129 10
rect -163 1 -129 4
rect -708 -2 -430 1
<< m2contact >>
rect -242 384 -237 389
rect -428 303 -423 308
rect -223 375 -218 380
rect -239 332 -234 337
rect -168 338 -163 343
rect -447 294 -442 299
rect -502 257 -497 262
rect -336 243 -331 248
rect -544 204 -539 209
rect -440 198 -435 203
rect -126 285 -121 290
rect -375 208 -370 213
rect -389 174 -384 179
rect -720 110 -715 115
rect -706 87 -701 92
rect -678 95 -673 100
rect -510 147 -505 152
rect -526 122 -521 127
rect -606 101 -601 106
rect -512 99 -507 104
rect -484 107 -479 112
rect -375 151 -370 156
rect -347 159 -342 164
rect -351 111 -346 116
rect -585 88 -580 93
rect -698 73 -693 78
rect -660 73 -655 78
rect -632 70 -627 75
rect -399 83 -394 89
rect -234 106 -229 111
rect -251 93 -246 98
rect -500 73 -495 78
rect -674 50 -669 55
rect -652 47 -647 52
rect -472 70 -467 75
rect -593 62 -588 67
rect -625 47 -620 52
rect -591 50 -586 55
rect -514 50 -509 55
rect -492 47 -487 52
rect -433 62 -428 67
rect -465 47 -460 52
rect -431 50 -426 55
rect -351 76 -346 81
rect -323 73 -318 78
rect -365 53 -360 58
rect -343 50 -338 55
rect -316 50 -311 55
rect -282 53 -277 58
rect -190 128 -185 133
rect -166 132 -161 137
rect -208 117 -203 122
rect -5 193 0 198
rect -24 187 -19 192
rect 25 170 30 175
rect 36 165 41 170
rect 90 170 95 175
rect 10 128 15 133
rect -217 107 -212 112
rect -180 109 -175 114
rect -132 91 -127 96
rect -199 76 -194 81
rect -171 73 -166 78
rect -114 82 -109 87
rect -213 53 -208 58
rect -191 50 -186 55
rect -132 65 -127 70
rect -164 50 -159 55
rect -130 53 -125 58
rect -79 87 -74 92
rect -41 87 -36 92
rect -76 51 -71 56
rect -82 24 -77 29
<< metal2 >>
rect -208 403 -205 416
rect -237 385 -220 388
rect -223 380 -220 385
rect -739 114 -736 366
rect -552 126 -549 365
rect -411 323 -408 375
rect -230 339 -168 342
rect -445 304 -428 307
rect -445 299 -442 304
rect -237 301 -234 332
rect -356 296 -345 299
rect -356 279 -353 296
rect -321 298 -234 301
rect -438 276 -353 279
rect -438 261 -435 276
rect -497 258 -435 261
rect -543 243 -484 246
rect -543 209 -540 243
rect -438 203 -435 258
rect -429 208 -426 257
rect -335 216 -332 243
rect -374 213 -332 216
rect -429 205 -416 208
rect -435 198 -424 201
rect -427 172 -424 198
rect -470 169 -424 172
rect -511 147 -510 150
rect -505 147 -501 150
rect -504 143 -501 147
rect -552 123 -526 126
rect -739 111 -720 114
rect -735 75 -732 102
rect -704 85 -701 87
rect -677 85 -674 95
rect -704 82 -674 85
rect -640 85 -637 119
rect -601 102 -585 105
rect -588 89 -585 102
rect -510 97 -507 99
rect -483 97 -480 107
rect -510 94 -480 97
rect -470 88 -467 169
rect -419 165 -416 205
rect -411 178 -407 211
rect -321 207 -318 298
rect -230 284 -227 339
rect -181 324 -122 327
rect -125 290 -122 324
rect -338 204 -318 207
rect -120 235 -16 238
rect -411 175 -389 178
rect -463 162 -416 165
rect -463 96 -460 162
rect -404 156 -401 166
rect -453 153 -401 156
rect -453 104 -450 153
rect -373 149 -370 151
rect -346 149 -343 159
rect -373 146 -343 149
rect -338 141 -335 204
rect -439 138 -335 141
rect -439 116 -436 138
rect -217 128 -190 131
rect -135 136 -132 178
rect -161 133 -132 136
rect -217 121 -214 128
rect -242 118 -214 121
rect -439 113 -374 116
rect -453 101 -385 104
rect -463 93 -395 96
rect -398 89 -395 93
rect -470 85 -429 88
rect -640 82 -589 85
rect -735 72 -709 75
rect -655 73 -632 74
rect -712 28 -709 72
rect -697 54 -694 73
rect -659 71 -632 73
rect -592 67 -589 82
rect -697 51 -674 54
rect -624 54 -621 56
rect -624 52 -591 54
rect -647 48 -625 51
rect -620 51 -591 52
rect -537 54 -534 74
rect -495 73 -472 74
rect -499 71 -472 73
rect -432 67 -429 85
rect -388 57 -385 101
rect -377 101 -374 113
rect -346 112 -315 115
rect -377 98 -326 101
rect -242 100 -239 118
rect -120 121 -117 235
rect -19 199 -16 235
rect -19 196 -12 199
rect -15 187 -12 196
rect -5 187 -2 193
rect -23 176 -20 187
rect -15 184 -2 187
rect -23 175 30 176
rect -23 173 25 175
rect 36 171 90 174
rect 36 170 41 171
rect -87 127 -76 130
rect -131 118 -117 121
rect -229 108 -217 111
rect -207 107 -204 117
rect -180 107 -177 109
rect -207 104 -177 107
rect -329 97 -326 98
rect -329 94 -251 97
rect -242 97 -233 100
rect -346 76 -323 77
rect -350 74 -323 76
rect -537 51 -514 54
rect -464 54 -461 56
rect -464 52 -431 54
rect -487 48 -465 51
rect -460 51 -431 52
rect -388 54 -365 57
rect -315 57 -312 59
rect -315 55 -282 57
rect -338 51 -316 54
rect -311 54 -282 55
rect -236 57 -233 97
rect -131 96 -128 118
rect -194 76 -171 77
rect -198 74 -171 76
rect -131 70 -128 91
rect -79 92 -76 127
rect -40 129 10 132
rect -40 92 -37 129
rect -109 83 -91 86
rect -236 54 -213 57
rect -163 57 -160 59
rect -163 55 -130 57
rect -186 51 -164 54
rect -159 54 -130 55
rect -94 55 -91 83
rect -94 52 -76 55
rect -712 25 -82 28
<< m3contact >>
rect -484 242 -479 247
rect -186 323 -181 328
rect -315 111 -310 116
rect -92 126 -87 131
<< m123contact >>
rect -561 259 -556 264
rect -665 146 -660 151
rect -141 348 -136 353
rect -159 343 -154 348
rect -333 323 -328 328
rect -283 319 -278 324
rect -529 267 -524 272
rect -490 203 -485 208
rect -430 257 -425 262
rect -387 238 -382 243
rect -439 187 -434 192
rect -528 175 -523 180
rect -640 119 -635 124
rect -736 102 -731 107
rect -705 104 -700 109
rect -590 116 -585 121
rect -542 114 -537 119
rect -511 116 -506 121
rect -559 104 -554 109
rect -230 279 -225 284
rect -186 279 -181 284
rect -231 270 -226 275
rect -142 256 -137 261
rect -123 248 -118 253
rect -405 166 -400 171
rect -374 168 -369 173
rect -145 164 -140 169
rect -234 136 -229 141
rect -181 126 -176 131
rect -150 124 -145 129
rect -690 58 -685 63
rect -625 61 -620 66
rect -659 56 -654 61
rect -559 56 -554 61
rect -530 58 -525 63
rect -465 61 -460 66
rect -499 56 -494 61
rect -5 202 0 207
rect 47 188 52 193
rect -29 163 -24 168
rect -381 61 -376 66
rect -316 64 -311 69
rect -284 65 -279 70
rect -350 59 -345 64
rect -99 90 -94 95
rect -229 61 -224 66
rect -164 64 -159 69
rect -198 59 -193 64
rect -250 52 -245 57
rect -591 35 -586 40
rect -431 35 -426 40
rect -282 38 -277 43
rect -130 38 -125 43
<< metal3 >>
rect -348 343 -159 346
rect -348 314 -345 343
rect -187 328 -180 329
rect -187 327 -186 328
rect -279 324 -186 327
rect -429 311 -345 314
rect -332 312 -329 323
rect -278 321 -276 324
rect -187 323 -186 324
rect -181 323 -180 328
rect -187 322 -180 323
rect -664 199 -609 202
rect -664 151 -661 199
rect -612 198 -609 199
rect -612 195 -588 198
rect -640 190 -624 193
rect -704 147 -665 150
rect -704 109 -701 147
rect -640 124 -637 190
rect -559 171 -556 259
rect -528 180 -525 267
rect -429 262 -426 311
rect -315 292 -240 295
rect -485 247 -478 248
rect -485 242 -484 247
rect -479 246 -478 247
rect -479 243 -386 246
rect -479 242 -478 243
rect -485 241 -478 242
rect -389 240 -387 243
rect -485 203 -483 208
rect -486 190 -483 203
rect -315 200 -312 292
rect -302 209 -299 292
rect -243 283 -240 292
rect -243 280 -230 283
rect -247 272 -231 275
rect -185 253 -182 279
rect -140 261 -137 348
rect -249 250 -182 253
rect -302 206 -222 209
rect -332 197 -312 200
rect -486 187 -475 190
rect -483 186 -480 187
rect -589 168 -556 171
rect -589 121 -586 168
rect -439 170 -435 187
rect -403 171 -374 172
rect -511 166 -435 170
rect -400 169 -374 171
rect -332 135 -329 197
rect -225 140 -222 206
rect -122 195 -119 248
rect -11 202 -5 206
rect -122 192 -108 195
rect -111 186 -108 192
rect -111 183 -72 186
rect -149 173 -142 176
rect -145 169 -142 173
rect -124 175 -83 178
rect -229 137 -222 140
rect -431 132 -329 135
rect -431 122 -428 132
rect -176 129 -147 130
rect -176 127 -150 129
rect -124 126 -121 175
rect -135 123 -121 126
rect -116 170 -108 171
rect -540 119 -511 120
rect -734 107 -705 108
rect -731 105 -705 107
rect -662 61 -625 64
rect -589 61 -586 116
rect -537 117 -511 119
rect -431 119 -367 122
rect -370 109 -367 119
rect -310 112 -304 115
rect -554 104 -550 108
rect -370 106 -319 109
rect -553 103 -550 104
rect -322 103 -319 106
rect -135 104 -132 123
rect -116 114 -113 170
rect -86 167 -83 175
rect -75 175 -72 183
rect -75 172 -25 175
rect -28 168 -25 172
rect -11 171 -8 202
rect -86 164 -35 167
rect -38 159 -35 164
rect 47 159 50 188
rect -38 156 50 159
rect -98 127 -92 130
rect -116 111 -106 114
rect -109 104 -106 111
rect -553 100 -552 103
rect -322 100 -280 103
rect -135 101 -115 104
rect -109 101 -86 104
rect -283 70 -280 100
rect -118 94 -115 101
rect -118 91 -99 94
rect -662 60 -659 61
rect -685 58 -659 60
rect -688 57 -659 58
rect -624 39 -621 61
rect -589 58 -559 61
rect -502 61 -465 64
rect -353 64 -316 67
rect -353 63 -350 64
rect -376 61 -350 63
rect -502 60 -499 61
rect -525 58 -499 60
rect -528 57 -499 58
rect -624 36 -591 39
rect -464 39 -461 61
rect -379 60 -350 61
rect -315 42 -312 64
rect -201 64 -164 67
rect -201 63 -198 64
rect -224 61 -198 63
rect -227 60 -198 61
rect -464 36 -431 39
rect -315 39 -282 42
rect -249 19 -246 52
rect -163 42 -160 64
rect -163 39 -130 42
rect -89 19 -86 101
rect -249 16 -86 19
<< m234contact >>
rect -209 398 -204 403
rect -412 318 -407 323
rect -345 295 -340 300
rect -412 211 -407 216
rect -516 166 -511 171
rect -505 138 -500 143
rect -136 178 -131 183
rect -538 74 -533 79
<< m4contact >>
rect -588 194 -583 199
rect -624 189 -619 194
rect -252 272 -247 277
rect -480 182 -475 187
rect -304 111 -299 116
rect -113 165 -108 170
rect -12 166 -7 171
rect -103 126 -98 131
<< metal4 >>
rect -411 216 -408 318
rect -340 295 -335 299
rect -338 289 -335 295
rect -338 286 -252 289
rect -255 272 -252 286
rect -583 196 -487 199
rect -619 190 -595 193
rect -598 170 -595 190
rect -490 185 -487 196
rect -208 190 -205 398
rect -208 187 -132 190
rect -490 182 -480 185
rect -135 183 -132 187
rect -598 167 -516 170
rect -108 166 -12 169
rect -504 87 -501 138
rect -111 126 -103 129
rect -111 119 -108 126
rect -111 116 -100 119
rect -299 112 -287 115
rect -290 107 -287 112
rect -103 107 -100 116
rect -290 104 -100 107
rect -537 84 -501 87
rect -537 79 -534 84
<< m345contact >>
rect -333 307 -328 312
rect -254 249 -249 254
rect -154 171 -149 176
rect -552 98 -547 103
<< metal5 >>
rect -332 294 -329 307
rect -332 291 -239 294
rect -309 281 -257 284
rect -309 210 -306 281
rect -299 274 -264 277
rect -299 213 -296 274
rect -267 244 -264 274
rect -260 254 -257 281
rect -260 250 -254 254
rect -242 244 -239 291
rect -267 241 -239 244
rect -299 210 -212 213
rect -336 207 -306 210
rect -336 164 -333 207
rect -215 175 -212 210
rect -215 172 -154 175
rect -468 161 -333 164
rect -468 102 -465 161
rect -547 99 -465 102
<< labels >>
rlabel metal1 -665 77 -665 77 1 b0_inv
rlabel metal1 -562 50 -556 53 7 g0_inv
rlabel metal1 -596 61 -592 64 1 p0_inv
rlabel metal1 -659 15 -657 18 1 b0
rlabel metal2 -697 75 -695 77 3 mid_s0
rlabel metal1 -684 56 -682 58 1 a0
rlabel metal1 -617 -1 -617 0 1 vdd
rlabel metal1 -607 81 -607 81 5 gnd
rlabel metal1 -687 87 -687 87 1 gnd
rlabel metal1 -718 108 -716 110 1 s0
rlabel metal1 -730 107 -728 109 1 c0
rlabel metal1 -697 106 -694 108 1 mid_s0
rlabel metal1 -562 119 -556 122 7 c1
rlabel metal1 -589 119 -585 121 1 g0_inv
rlabel metal1 -569 90 -569 90 1 gnd
rlabel metal1 -595 126 -593 129 1 temp100
rlabel metal1 -622 104 -622 104 1 gnd
rlabel metal1 -647 148 -645 151 1 c0_inv
rlabel metal1 -662 147 -660 149 3 c0
rlabel metal1 -472 19 -472 19 1 vdd
rlabel metal1 -447 81 -447 81 5 gnd
rlabel metal1 -457 -1 -457 0 1 vdd
rlabel metal1 -418 9 -418 9 1 vdd
rlabel metal2 -537 75 -535 77 3 mid_s1
rlabel metal1 -524 56 -522 58 1 a1
rlabel metal1 -499 15 -497 18 1 b1
rlabel metal1 -436 61 -432 64 1 p1_inv
rlabel metal1 -402 50 -396 53 7 g1_inv
rlabel m2contact -498 76 -496 78 1 b1_inv
rlabel metal1 -524 120 -522 122 1 s1
rlabel metal1 -484 158 -484 158 5 vdd
rlabel metal1 -443 256 -443 257 5 vdd
rlabel metal1 -453 175 -453 175 1 gnd
rlabel metal1 -442 198 -438 200 7 p1_inv
rlabel metal1 -441 192 -436 194 7 p0_inv
rlabel metal1 -469 196 -465 198 3 temp101
rlabel metal1 -499 250 -499 250 5 vdd
rlabel metal1 -508 177 -508 177 1 gnd
rlabel metal1 -492 206 -488 207 1 c0
rlabel metal1 -536 207 -534 209 1 temp102
rlabel metal1 -525 279 -525 279 3 gnd
rlabel metal1 -444 269 -443 269 7 vdd
rlabel metal1 -503 305 -500 308 1 temp103
rlabel metal1 -416 304 -416 304 5 vdd
rlabel metal1 -407 231 -407 231 1 gnd
rlabel metal1 -424 260 -424 260 1 g1_inv
rlabel metal1 -400 260 -394 263 7 temp104
rlabel metal1 -378 304 -378 305 5 vdd
rlabel metal1 -368 223 -368 223 1 gnd
rlabel metal1 -341 245 -339 247 1 c2
rlabel metal1 -508 261 -505 264 1 g0_inv
rlabel metal1 -639 121 -634 124 1 p0_inv
rlabel metal1 -350 18 -348 21 1 b2
rlabel metal1 -375 59 -373 61 1 a2
rlabel metal2 -388 78 -386 80 3 mid_s2
rlabel m2contact -349 79 -347 81 1 b2_inv
rlabel metal1 -287 64 -283 67 1 p2_inv
rlabel metal1 -253 53 -247 56 7 g2_inv
rlabel metal1 -269 12 -269 12 1 vdd
rlabel metal1 -308 2 -308 3 1 vdd
rlabel metal1 -298 84 -298 84 5 gnd
rlabel metal1 -323 22 -323 22 1 vdd
rlabel metal1 -387 172 -385 174 1 s2
rlabel metal1 -356 151 -356 151 1 gnd
rlabel metal1 -222 337 -222 338 5 vdd
rlabel metal1 -212 256 -212 256 1 gnd
rlabel metal1 -166 331 -166 331 5 vdd
rlabel metal1 -157 258 -157 258 1 gnd
rlabel metal1 -140 360 -140 360 7 gnd
rlabel metal1 -222 350 -221 350 3 vdd
rlabel metal1 -249 385 -249 385 5 vdd
rlabel metal1 -258 312 -258 312 1 gnd
rlabel metal1 -287 385 -287 386 5 vdd
rlabel metal1 -297 304 -297 304 1 gnd
rlabel metal1 -326 326 -324 328 1 c3
rlabel metal1 -271 341 -265 344 1 temp108
rlabel metal1 -131 288 -129 290 1 temp106
rlabel metal1 -177 287 -173 288 1 c1
rlabel metal1 -200 277 -196 279 1 temp105
rlabel metal1 -227 279 -223 281 1 p2_inv
rlabel metal1 -165 386 -162 389 1 temp107
rlabel metal1 -242 340 -240 342 1 g2_inv
rlabel metal1 -159 344 -156 347 1 g1_inv
rlabel metal1 -225 274 -225 274 1 p1_inv
rlabel metal1 -236 202 -236 203 5 vdd
rlabel metal1 -246 121 -246 121 1 gnd
rlabel metal1 -235 144 -231 146 7 p3_inv
rlabel metal1 -261 142 -260 144 3 temp109
rlabel metal1 -278 197 -278 197 5 vdd
rlabel metal1 -287 124 -287 124 1 gnd
rlabel metal1 -271 159 -268 162 1 temp101
rlabel metal1 -315 154 -313 156 1 p4
rlabel metal1 -171 22 -171 22 1 vdd
rlabel metal1 -146 84 -146 84 5 gnd
rlabel metal1 -156 2 -156 3 1 vdd
rlabel metal1 -117 12 -117 12 1 vdd
rlabel m2contact -197 79 -195 81 1 b3_inv
rlabel metal2 -236 78 -234 80 3 mid_s3
rlabel metal1 -223 59 -221 61 1 a3
rlabel metal1 -198 18 -196 21 1 b3
rlabel metal1 -101 53 -95 56 7 g3_inv
rlabel metal1 -135 64 -131 67 1 p3_inv
rlabel m123contact -232 139 -232 139 1 p2_inv
rlabel metal1 -358 208 -358 208 1 vdd
rlabel metal3 -152 130 -152 130 1 in2
rlabel metal1 -194 109 -194 109 1 gnd
rlabel metal1 -203 168 -203 168 5 vdd
rlabel metal1 -165 130 -163 132 1 s3
rlabel metal1 33 134 35 137 1 g4_inv
rlabel metal1 56 150 56 150 7 gnd
rlabel metal1 -26 160 -25 160 3 vdd
rlabel metal1 83 195 89 198 7 temp112
rlabel metal1 57 194 59 197 1 g3_inv
rlabel metal1 76 166 76 166 1 gnd
rlabel metal1 67 239 67 239 5 vdd
rlabel m2contact -1 196 -1 196 1 p3_inv
rlabel metal1 40 202 42 204 1 temp111
rlabel metal1 13 180 13 180 1 gnd
rlabel metal1 3 261 3 262 5 vdd
rlabel metal1 -116 212 -116 212 1 temp110
rlabel metal1 -76 213 -64 216 1 temp104
rlabel metal1 -70 208 -70 208 1 temp109
rlabel metal1 -77 271 -77 272 5 vdd
rlabel metal1 -87 190 -87 190 1 gnd
rlabel metal1 -22 208 -22 210 1 temp110
rlabel metal1 -49 178 -49 178 1 gnd
rlabel metal1 -58 251 -58 251 5 vdd
rlabel metal1 -63 126 -63 126 5 vdd
rlabel metal1 -54 53 -54 53 1 gnd
rlabel metal1 -72 88 -70 91 3 p4
rlabel metal1 -73 81 -70 84 3 c0
rlabel metal1 -29 126 -29 126 5 vdd
rlabel metal1 -20 53 -20 53 1 gnd
rlabel metal1 -37 82 -35 83 1 temp113
rlabel m2contact -39 88 -36 91 1 g4_inv
rlabel metal1 -13 82 -7 85 7 c4
<< end >>
